localparam NUM_PIXELS_TARGET6 = 16;
logic [23:0] target6 [0:15];
assign target6[0] = 24'hffff00;
assign target6[1] = 24'hffff00;
assign target6[2] = 24'h000000;
assign target6[3] = 24'h000000;
assign target6[4] = 24'hffff00;
assign target6[5] = 24'hffff00;
assign target6[6] = 24'h000000;
assign target6[7] = 24'h000000;
assign target6[8] = 24'hffff00;
assign target6[9] = 24'hffff00;
assign target6[10] = 24'h000000;
assign target6[11] = 24'h000000;
assign target6[12] = 24'hffff00;
assign target6[13] = 24'hffff00;
assign target6[14] = 24'h000000;
assign target6[15] = 24'h000000;
