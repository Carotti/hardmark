localparam NUM_PIXELS_TARGET1 = 16;
logic [23:0] target1 [0:15];
assign target1[0] = 24'h000000;
assign target1[1] = 24'h000000;
assign target1[2] = 24'h000000;
assign target1[3] = 24'h000000;
assign target1[4] = 24'hffffff;
assign target1[5] = 24'hffffff;
assign target1[6] = 24'hffffff;
assign target1[7] = 24'hffffff;
assign target1[8] = 24'h000000;
assign target1[9] = 24'h000000;
assign target1[10] = 24'h000000;
assign target1[11] = 24'h000000;
assign target1[12] = 24'hffffff;
assign target1[13] = 24'hffffff;
assign target1[14] = 24'hffffff;
assign target1[15] = 24'hffffff;
