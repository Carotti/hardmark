`include "target2.sv"
`include "full_test1.sv"
`include "target6.sv"
`include "target3.sv"
`include "target_only_stripe.sv"
`include "target1.sv"
`include "target7.sv"
`include "target4.sv"
`include "target5.sv"
