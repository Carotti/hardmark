localparam NUM_PIXELS_TARGET3 = 16;
logic [23:0] target3 [0:15];
assign target3[0] = 24'h000000;
assign target3[1] = 24'hffffff;
assign target3[2] = 24'hffffff;
assign target3[3] = 24'hffffff;
assign target3[4] = 24'hffffff;
assign target3[5] = 24'h000000;
assign target3[6] = 24'hffffff;
assign target3[7] = 24'hffffff;
assign target3[8] = 24'hffffff;
assign target3[9] = 24'hffffff;
assign target3[10] = 24'h000000;
assign target3[11] = 24'hffffff;
assign target3[12] = 24'hffffff;
assign target3[13] = 24'hffffff;
assign target3[14] = 24'hffffff;
assign target3[15] = 24'h000000;
