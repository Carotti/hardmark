`include "full_test1.sv"
