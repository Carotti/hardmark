localparam NUM_PIXELS_TARGET4 = 16;
logic [23:0] target4 [0:15];
assign target4[0] = 24'h00ffff;
assign target4[1] = 24'h00ffff;
assign target4[2] = 24'h000000;
assign target4[3] = 24'h000000;
assign target4[4] = 24'h00ffff;
assign target4[5] = 24'h00ffff;
assign target4[6] = 24'h000000;
assign target4[7] = 24'h000000;
assign target4[8] = 24'h00ffff;
assign target4[9] = 24'h00ffff;
assign target4[10] = 24'h000000;
assign target4[11] = 24'h000000;
assign target4[12] = 24'h00ffff;
assign target4[13] = 24'h00ffff;
assign target4[14] = 24'h000000;
assign target4[15] = 24'h000000;
