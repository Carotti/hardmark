localparam NUM_PIXELS_TARGET2 = 16;
logic [23:0] target2 [0:15];
assign target2[0] = 24'h000000;
assign target2[1] = 24'hffffff;
assign target2[2] = 24'h000000;
assign target2[3] = 24'hffffff;
assign target2[4] = 24'h000000;
assign target2[5] = 24'hffffff;
assign target2[6] = 24'h000000;
assign target2[7] = 24'hffffff;
assign target2[8] = 24'h000000;
assign target2[9] = 24'hffffff;
assign target2[10] = 24'h000000;
assign target2[11] = 24'hffffff;
assign target2[12] = 24'h000000;
assign target2[13] = 24'hffffff;
assign target2[14] = 24'h000000;
assign target2[15] = 24'hffffff;
