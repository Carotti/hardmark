localparam NUM_PIXELS_TARGET5 = 16;
logic [23:0] target5 [0:15];
assign target5[0] = 24'hff00ff;
assign target5[1] = 24'hff00ff;
assign target5[2] = 24'h000000;
assign target5[3] = 24'h000000;
assign target5[4] = 24'hff00ff;
assign target5[5] = 24'hff00ff;
assign target5[6] = 24'h000000;
assign target5[7] = 24'h000000;
assign target5[8] = 24'hff00ff;
assign target5[9] = 24'hff00ff;
assign target5[10] = 24'h000000;
assign target5[11] = 24'h000000;
assign target5[12] = 24'hff00ff;
assign target5[13] = 24'hff00ff;
assign target5[14] = 24'h000000;
assign target5[15] = 24'h000000;
