localparam NUM_PIXELS_TARGET_ONLY_STRIPE = 9212;
logic [23:0] target_only_stripe [0:9211];
assign target_only_stripe[0] = 24'h000000;
assign target_only_stripe[1] = 24'h000000;
assign target_only_stripe[2] = 24'h000000;
assign target_only_stripe[3] = 24'h000000;
assign target_only_stripe[4] = 24'h000000;
assign target_only_stripe[5] = 24'h000000;
assign target_only_stripe[6] = 24'h000000;
assign target_only_stripe[7] = 24'h000000;
assign target_only_stripe[8] = 24'h000000;
assign target_only_stripe[9] = 24'h000000;
assign target_only_stripe[10] = 24'h000000;
assign target_only_stripe[11] = 24'h000000;
assign target_only_stripe[12] = 24'h000000;
assign target_only_stripe[13] = 24'h000000;
assign target_only_stripe[14] = 24'h000000;
assign target_only_stripe[15] = 24'h000000;
assign target_only_stripe[16] = 24'h000000;
assign target_only_stripe[17] = 24'h000000;
assign target_only_stripe[18] = 24'h000000;
assign target_only_stripe[19] = 24'h000000;
assign target_only_stripe[20] = 24'h000000;
assign target_only_stripe[21] = 24'h000000;
assign target_only_stripe[22] = 24'h000000;
assign target_only_stripe[23] = 24'h000000;
assign target_only_stripe[24] = 24'h000000;
assign target_only_stripe[25] = 24'h000000;
assign target_only_stripe[26] = 24'h000000;
assign target_only_stripe[27] = 24'h000000;
assign target_only_stripe[28] = 24'h000000;
assign target_only_stripe[29] = 24'h000000;
assign target_only_stripe[30] = 24'h000000;
assign target_only_stripe[31] = 24'h000000;
assign target_only_stripe[32] = 24'ha5a5a5;
assign target_only_stripe[33] = 24'hffffff;
assign target_only_stripe[34] = 24'hffffff;
assign target_only_stripe[35] = 24'hffffff;
assign target_only_stripe[36] = 24'hffffff;
assign target_only_stripe[37] = 24'hffffff;
assign target_only_stripe[38] = 24'hffffff;
assign target_only_stripe[39] = 24'hffffff;
assign target_only_stripe[40] = 24'hffffff;
assign target_only_stripe[41] = 24'hffffff;
assign target_only_stripe[42] = 24'hffffff;
assign target_only_stripe[43] = 24'hffffff;
assign target_only_stripe[44] = 24'hffffff;
assign target_only_stripe[45] = 24'hffffff;
assign target_only_stripe[46] = 24'hffffff;
assign target_only_stripe[47] = 24'hffffff;
assign target_only_stripe[48] = 24'hffffff;
assign target_only_stripe[49] = 24'hffffff;
assign target_only_stripe[50] = 24'hffffff;
assign target_only_stripe[51] = 24'hffffff;
assign target_only_stripe[52] = 24'hffffff;
assign target_only_stripe[53] = 24'hfaf7f5;
assign target_only_stripe[54] = 24'hebe6db;
assign target_only_stripe[55] = 24'hebe6db;
assign target_only_stripe[56] = 24'hfaf9f7;
assign target_only_stripe[57] = 24'hffffff;
assign target_only_stripe[58] = 24'hffffff;
assign target_only_stripe[59] = 24'hffffff;
assign target_only_stripe[60] = 24'hffffff;
assign target_only_stripe[61] = 24'hffffff;
assign target_only_stripe[62] = 24'hffffff;
assign target_only_stripe[63] = 24'hffffff;
assign target_only_stripe[64] = 24'hffffff;
assign target_only_stripe[65] = 24'hffffff;
assign target_only_stripe[66] = 24'hffffff;
assign target_only_stripe[67] = 24'h000000;
assign target_only_stripe[68] = 24'h000000;
assign target_only_stripe[69] = 24'h000000;
assign target_only_stripe[70] = 24'h000000;
assign target_only_stripe[71] = 24'h000000;
assign target_only_stripe[72] = 24'h000000;
assign target_only_stripe[73] = 24'h000000;
assign target_only_stripe[74] = 24'h000000;
assign target_only_stripe[75] = 24'h000000;
assign target_only_stripe[76] = 24'h000000;
assign target_only_stripe[77] = 24'h000000;
assign target_only_stripe[78] = 24'h000000;
assign target_only_stripe[79] = 24'h000000;
assign target_only_stripe[80] = 24'h000000;
assign target_only_stripe[81] = 24'h000000;
assign target_only_stripe[82] = 24'h000000;
assign target_only_stripe[83] = 24'h000000;
assign target_only_stripe[84] = 24'h000000;
assign target_only_stripe[85] = 24'h000000;
assign target_only_stripe[86] = 24'h000000;
assign target_only_stripe[87] = 24'h000000;
assign target_only_stripe[88] = 24'h000000;
assign target_only_stripe[89] = 24'h000000;
assign target_only_stripe[90] = 24'h000000;
assign target_only_stripe[91] = 24'h000000;
assign target_only_stripe[92] = 24'h000000;
assign target_only_stripe[93] = 24'h000000;
assign target_only_stripe[94] = 24'h000000;
assign target_only_stripe[95] = 24'h000000;
assign target_only_stripe[96] = 24'h000000;
assign target_only_stripe[97] = 24'h000000;
assign target_only_stripe[98] = 24'h000000;
assign target_only_stripe[99] = 24'haeaeae;
assign target_only_stripe[100] = 24'hffffff;
assign target_only_stripe[101] = 24'hffffff;
assign target_only_stripe[102] = 24'hffffff;
assign target_only_stripe[103] = 24'hffffff;
assign target_only_stripe[104] = 24'hffffff;
assign target_only_stripe[105] = 24'hffffff;
assign target_only_stripe[106] = 24'hffffff;
assign target_only_stripe[107] = 24'hffffff;
assign target_only_stripe[108] = 24'hffffff;
assign target_only_stripe[109] = 24'hffffff;
assign target_only_stripe[110] = 24'hffffff;
assign target_only_stripe[111] = 24'hffffff;
assign target_only_stripe[112] = 24'hffffff;
assign target_only_stripe[113] = 24'hffffff;
assign target_only_stripe[114] = 24'hffffff;
assign target_only_stripe[115] = 24'hffffff;
assign target_only_stripe[116] = 24'hffffff;
assign target_only_stripe[117] = 24'hffffff;
assign target_only_stripe[118] = 24'hffffff;
assign target_only_stripe[119] = 24'hffffff;
assign target_only_stripe[120] = 24'hffffff;
assign target_only_stripe[121] = 24'hffffff;
assign target_only_stripe[122] = 24'hffffff;
assign target_only_stripe[123] = 24'hffffff;
assign target_only_stripe[124] = 24'hffffff;
assign target_only_stripe[125] = 24'hffffff;
assign target_only_stripe[126] = 24'hffffff;
assign target_only_stripe[127] = 24'hffffff;
assign target_only_stripe[128] = 24'hffffff;
assign target_only_stripe[129] = 24'hffffff;
assign target_only_stripe[130] = 24'hffffff;
assign target_only_stripe[131] = 24'hffffff;
assign target_only_stripe[132] = 24'hffffff;
assign target_only_stripe[133] = 24'hffffff;
assign target_only_stripe[134] = 24'hffffff;
assign target_only_stripe[135] = 24'h000000;
assign target_only_stripe[136] = 24'h000000;
assign target_only_stripe[137] = 24'h000000;
assign target_only_stripe[138] = 24'h000000;
assign target_only_stripe[139] = 24'h000000;
assign target_only_stripe[140] = 24'h000000;
assign target_only_stripe[141] = 24'h000000;
assign target_only_stripe[142] = 24'h000000;
assign target_only_stripe[143] = 24'h000000;
assign target_only_stripe[144] = 24'h000000;
assign target_only_stripe[145] = 24'h000000;
assign target_only_stripe[146] = 24'h000000;
assign target_only_stripe[147] = 24'h000000;
assign target_only_stripe[148] = 24'h000000;
assign target_only_stripe[149] = 24'h000000;
assign target_only_stripe[150] = 24'h000000;
assign target_only_stripe[151] = 24'h000000;
assign target_only_stripe[152] = 24'h000000;
assign target_only_stripe[153] = 24'h000000;
assign target_only_stripe[154] = 24'h000000;
assign target_only_stripe[155] = 24'h000000;
assign target_only_stripe[156] = 24'h000000;
assign target_only_stripe[157] = 24'h000000;
assign target_only_stripe[158] = 24'h000000;
assign target_only_stripe[159] = 24'h000000;
assign target_only_stripe[160] = 24'h000000;
assign target_only_stripe[161] = 24'h000000;
assign target_only_stripe[162] = 24'h000000;
assign target_only_stripe[163] = 24'h000000;
assign target_only_stripe[164] = 24'h000000;
assign target_only_stripe[165] = 24'h000000;
assign target_only_stripe[166] = 24'h000000;
assign target_only_stripe[167] = 24'h000000;
assign target_only_stripe[168] = 24'h000000;
assign target_only_stripe[169] = 24'h000000;
assign target_only_stripe[170] = 24'h000000;
assign target_only_stripe[171] = 24'h000000;
assign target_only_stripe[172] = 24'h000000;
assign target_only_stripe[173] = 24'h000000;
assign target_only_stripe[174] = 24'h000000;
assign target_only_stripe[175] = 24'h000000;
assign target_only_stripe[176] = 24'h000000;
assign target_only_stripe[177] = 24'h000000;
assign target_only_stripe[178] = 24'h000000;
assign target_only_stripe[179] = 24'h000000;
assign target_only_stripe[180] = 24'h000000;
assign target_only_stripe[181] = 24'h000000;
assign target_only_stripe[182] = 24'h000000;
assign target_only_stripe[183] = 24'h000000;
assign target_only_stripe[184] = 24'h000000;
assign target_only_stripe[185] = 24'h000000;
assign target_only_stripe[186] = 24'h000000;
assign target_only_stripe[187] = 24'h000000;
assign target_only_stripe[188] = 24'h000000;
assign target_only_stripe[189] = 24'h000000;
assign target_only_stripe[190] = 24'h000000;
assign target_only_stripe[191] = 24'h000000;
assign target_only_stripe[192] = 24'h000000;
assign target_only_stripe[193] = 24'h000000;
assign target_only_stripe[194] = 24'h818181;
assign target_only_stripe[195] = 24'hffffff;
assign target_only_stripe[196] = 24'hffffff;
assign target_only_stripe[197] = 24'hffffff;
assign target_only_stripe[198] = 24'hffffff;
assign target_only_stripe[199] = 24'hffffff;
assign target_only_stripe[200] = 24'hffffff;
assign target_only_stripe[201] = 24'hffffff;
assign target_only_stripe[202] = 24'hffffff;
assign target_only_stripe[203] = 24'hffffff;
assign target_only_stripe[204] = 24'hffffff;
assign target_only_stripe[205] = 24'hffffff;
assign target_only_stripe[206] = 24'hffffff;
assign target_only_stripe[207] = 24'hffffff;
assign target_only_stripe[208] = 24'hffffff;
assign target_only_stripe[209] = 24'hffffff;
assign target_only_stripe[210] = 24'hffffff;
assign target_only_stripe[211] = 24'hffffff;
assign target_only_stripe[212] = 24'hffffff;
assign target_only_stripe[213] = 24'hffffff;
assign target_only_stripe[214] = 24'hffffff;
assign target_only_stripe[215] = 24'hffffff;
assign target_only_stripe[216] = 24'hffffff;
assign target_only_stripe[217] = 24'hffffff;
assign target_only_stripe[218] = 24'hffffff;
assign target_only_stripe[219] = 24'hffffff;
assign target_only_stripe[220] = 24'hffffff;
assign target_only_stripe[221] = 24'hffffff;
assign target_only_stripe[222] = 24'hffffff;
assign target_only_stripe[223] = 24'hffffff;
assign target_only_stripe[224] = 24'hffffff;
assign target_only_stripe[225] = 24'hffffff;
assign target_only_stripe[226] = 24'hffffff;
assign target_only_stripe[227] = 24'hffffff;
assign target_only_stripe[228] = 24'hffffff;
assign target_only_stripe[229] = 24'hbdbdbd;
assign target_only_stripe[230] = 24'h000000;
assign target_only_stripe[231] = 24'h000000;
assign target_only_stripe[232] = 24'h000000;
assign target_only_stripe[233] = 24'h000000;
assign target_only_stripe[234] = 24'h000000;
assign target_only_stripe[235] = 24'h000000;
assign target_only_stripe[236] = 24'h000000;
assign target_only_stripe[237] = 24'h000000;
assign target_only_stripe[238] = 24'h000000;
assign target_only_stripe[239] = 24'h000000;
assign target_only_stripe[240] = 24'h000000;
assign target_only_stripe[241] = 24'h000000;
assign target_only_stripe[242] = 24'h000000;
assign target_only_stripe[243] = 24'h000000;
assign target_only_stripe[244] = 24'h000000;
assign target_only_stripe[245] = 24'h000000;
assign target_only_stripe[246] = 24'h000000;
assign target_only_stripe[247] = 24'h000000;
assign target_only_stripe[248] = 24'h000000;
assign target_only_stripe[249] = 24'h000000;
assign target_only_stripe[250] = 24'h000000;
assign target_only_stripe[251] = 24'h000000;
assign target_only_stripe[252] = 24'h000000;
assign target_only_stripe[253] = 24'h000000;
assign target_only_stripe[254] = 24'h000000;
assign target_only_stripe[255] = 24'h000000;
assign target_only_stripe[256] = 24'h000000;
assign target_only_stripe[257] = 24'h000000;
assign target_only_stripe[258] = 24'h000000;
assign target_only_stripe[259] = 24'h000000;
assign target_only_stripe[260] = 24'h000000;
assign target_only_stripe[261] = 24'h000000;
assign target_only_stripe[262] = 24'hffffff;
assign target_only_stripe[263] = 24'hffffff;
assign target_only_stripe[264] = 24'hffffff;
assign target_only_stripe[265] = 24'hfaf7f5;
assign target_only_stripe[266] = 24'hffffff;
assign target_only_stripe[267] = 24'hffffff;
assign target_only_stripe[268] = 24'hffffff;
assign target_only_stripe[269] = 24'hffffff;
assign target_only_stripe[270] = 24'hffffff;
assign target_only_stripe[271] = 24'hffffff;
assign target_only_stripe[272] = 24'hffffff;
assign target_only_stripe[273] = 24'hffffff;
assign target_only_stripe[274] = 24'hffffff;
assign target_only_stripe[275] = 24'hffffff;
assign target_only_stripe[276] = 24'hffffff;
assign target_only_stripe[277] = 24'hffffff;
assign target_only_stripe[278] = 24'hffffff;
assign target_only_stripe[279] = 24'hffffff;
assign target_only_stripe[280] = 24'hffffff;
assign target_only_stripe[281] = 24'hffffff;
assign target_only_stripe[282] = 24'hffffff;
assign target_only_stripe[283] = 24'hffffff;
assign target_only_stripe[284] = 24'hffffff;
assign target_only_stripe[285] = 24'hffffff;
assign target_only_stripe[286] = 24'hffffff;
assign target_only_stripe[287] = 24'hffffff;
assign target_only_stripe[288] = 24'hffffff;
assign target_only_stripe[289] = 24'hffffff;
assign target_only_stripe[290] = 24'hffffff;
assign target_only_stripe[291] = 24'hffffff;
assign target_only_stripe[292] = 24'hffffff;
assign target_only_stripe[293] = 24'hffffff;
assign target_only_stripe[294] = 24'hffffff;
assign target_only_stripe[295] = 24'hffffff;
assign target_only_stripe[296] = 24'hacacac;
assign target_only_stripe[297] = 24'h000000;
assign target_only_stripe[298] = 24'h000000;
assign target_only_stripe[299] = 24'h000000;
assign target_only_stripe[300] = 24'h000000;
assign target_only_stripe[301] = 24'h000000;
assign target_only_stripe[302] = 24'h000000;
assign target_only_stripe[303] = 24'h000000;
assign target_only_stripe[304] = 24'h000000;
assign target_only_stripe[305] = 24'h000000;
assign target_only_stripe[306] = 24'h000000;
assign target_only_stripe[307] = 24'h000000;
assign target_only_stripe[308] = 24'h000000;
assign target_only_stripe[309] = 24'h000000;
assign target_only_stripe[310] = 24'h000000;
assign target_only_stripe[311] = 24'h000000;
assign target_only_stripe[312] = 24'h000000;
assign target_only_stripe[313] = 24'h000000;
assign target_only_stripe[314] = 24'h000000;
assign target_only_stripe[315] = 24'h000000;
assign target_only_stripe[316] = 24'h000000;
assign target_only_stripe[317] = 24'h000000;
assign target_only_stripe[318] = 24'h000000;
assign target_only_stripe[319] = 24'h000000;
assign target_only_stripe[320] = 24'h000000;
assign target_only_stripe[321] = 24'h000000;
assign target_only_stripe[322] = 24'h000000;
assign target_only_stripe[323] = 24'h000000;
assign target_only_stripe[324] = 24'h000000;
assign target_only_stripe[325] = 24'h000000;
assign target_only_stripe[326] = 24'h000000;
assign target_only_stripe[327] = 24'h000000;
assign target_only_stripe[328] = 24'h000000;
assign target_only_stripe[329] = 24'h000000;
assign target_only_stripe[330] = 24'h000000;
assign target_only_stripe[331] = 24'h000000;
assign target_only_stripe[332] = 24'h000000;
assign target_only_stripe[333] = 24'h000000;
assign target_only_stripe[334] = 24'h000000;
assign target_only_stripe[335] = 24'h000000;
assign target_only_stripe[336] = 24'h000000;
assign target_only_stripe[337] = 24'h000000;
assign target_only_stripe[338] = 24'h000000;
assign target_only_stripe[339] = 24'h000000;
assign target_only_stripe[340] = 24'h000000;
assign target_only_stripe[341] = 24'h000000;
assign target_only_stripe[342] = 24'h000000;
assign target_only_stripe[343] = 24'h000000;
assign target_only_stripe[344] = 24'h000000;
assign target_only_stripe[345] = 24'h000000;
assign target_only_stripe[346] = 24'h000000;
assign target_only_stripe[347] = 24'h000000;
assign target_only_stripe[348] = 24'h000000;
assign target_only_stripe[349] = 24'h000000;
assign target_only_stripe[350] = 24'h000000;
assign target_only_stripe[351] = 24'h000000;
assign target_only_stripe[352] = 24'h000000;
assign target_only_stripe[353] = 24'h000000;
assign target_only_stripe[354] = 24'h000000;
assign target_only_stripe[355] = 24'h000000;
assign target_only_stripe[356] = 24'h000000;
assign target_only_stripe[357] = 24'h000000;
assign target_only_stripe[358] = 24'h000000;
assign target_only_stripe[359] = 24'h000000;
assign target_only_stripe[360] = 24'h000000;
assign target_only_stripe[361] = 24'hb2b2b2;
assign target_only_stripe[362] = 24'hffffff;
assign target_only_stripe[363] = 24'hffffff;
assign target_only_stripe[364] = 24'hffffff;
assign target_only_stripe[365] = 24'hffffff;
assign target_only_stripe[366] = 24'hffffff;
assign target_only_stripe[367] = 24'hffffff;
assign target_only_stripe[368] = 24'hffffff;
assign target_only_stripe[369] = 24'hffffff;
assign target_only_stripe[370] = 24'hffffff;
assign target_only_stripe[371] = 24'hffffff;
assign target_only_stripe[372] = 24'hffffff;
assign target_only_stripe[373] = 24'hffffff;
assign target_only_stripe[374] = 24'hffffff;
assign target_only_stripe[375] = 24'hffffff;
assign target_only_stripe[376] = 24'hffffff;
assign target_only_stripe[377] = 24'hffffff;
assign target_only_stripe[378] = 24'hffffff;
assign target_only_stripe[379] = 24'hffffff;
assign target_only_stripe[380] = 24'hffffff;
assign target_only_stripe[381] = 24'hffffff;
assign target_only_stripe[382] = 24'hffffff;
assign target_only_stripe[383] = 24'hede6db;
assign target_only_stripe[384] = 24'hf0e8de;
assign target_only_stripe[385] = 24'hede6db;
assign target_only_stripe[386] = 24'hffffff;
assign target_only_stripe[387] = 24'hffffff;
assign target_only_stripe[388] = 24'hffffff;
assign target_only_stripe[389] = 24'hffffff;
assign target_only_stripe[390] = 24'hffffff;
assign target_only_stripe[391] = 24'hffffff;
assign target_only_stripe[392] = 24'hffffff;
assign target_only_stripe[393] = 24'hffffff;
assign target_only_stripe[394] = 24'hffffff;
assign target_only_stripe[395] = 24'he7e7e7;
assign target_only_stripe[396] = 24'h000000;
assign target_only_stripe[397] = 24'h000000;
assign target_only_stripe[398] = 24'h000000;
assign target_only_stripe[399] = 24'h000000;
assign target_only_stripe[400] = 24'h000000;
assign target_only_stripe[401] = 24'h000000;
assign target_only_stripe[402] = 24'h000000;
assign target_only_stripe[403] = 24'h000000;
assign target_only_stripe[404] = 24'h000000;
assign target_only_stripe[405] = 24'h000000;
assign target_only_stripe[406] = 24'h000000;
assign target_only_stripe[407] = 24'h000000;
assign target_only_stripe[408] = 24'h000000;
assign target_only_stripe[409] = 24'h000000;
assign target_only_stripe[410] = 24'h000000;
assign target_only_stripe[411] = 24'h000000;
assign target_only_stripe[412] = 24'h000000;
assign target_only_stripe[413] = 24'h000000;
assign target_only_stripe[414] = 24'h000000;
assign target_only_stripe[415] = 24'h000000;
assign target_only_stripe[416] = 24'h000000;
assign target_only_stripe[417] = 24'h000000;
assign target_only_stripe[418] = 24'h000000;
assign target_only_stripe[419] = 24'h000000;
assign target_only_stripe[420] = 24'h000000;
assign target_only_stripe[421] = 24'h000000;
assign target_only_stripe[422] = 24'h000000;
assign target_only_stripe[423] = 24'h000000;
assign target_only_stripe[424] = 24'h000000;
assign target_only_stripe[425] = 24'h000000;
assign target_only_stripe[426] = 24'h000000;
assign target_only_stripe[427] = 24'h010101;
assign target_only_stripe[428] = 24'hfbfbfb;
assign target_only_stripe[429] = 24'hffffff;
assign target_only_stripe[430] = 24'hffffff;
assign target_only_stripe[431] = 24'hffffff;
assign target_only_stripe[432] = 24'hffffff;
assign target_only_stripe[433] = 24'hffffff;
assign target_only_stripe[434] = 24'hffffff;
assign target_only_stripe[435] = 24'hffffff;
assign target_only_stripe[436] = 24'hffffff;
assign target_only_stripe[437] = 24'hffffff;
assign target_only_stripe[438] = 24'hffffff;
assign target_only_stripe[439] = 24'hffffff;
assign target_only_stripe[440] = 24'hffffff;
assign target_only_stripe[441] = 24'hffffff;
assign target_only_stripe[442] = 24'hffffff;
assign target_only_stripe[443] = 24'hffffff;
assign target_only_stripe[444] = 24'hffffff;
assign target_only_stripe[445] = 24'hffffff;
assign target_only_stripe[446] = 24'hffffff;
assign target_only_stripe[447] = 24'hffffff;
assign target_only_stripe[448] = 24'hffffff;
assign target_only_stripe[449] = 24'hffffff;
assign target_only_stripe[450] = 24'hffffff;
assign target_only_stripe[451] = 24'hffffff;
assign target_only_stripe[452] = 24'hffffff;
assign target_only_stripe[453] = 24'hffffff;
assign target_only_stripe[454] = 24'hffffff;
assign target_only_stripe[455] = 24'hffffff;
assign target_only_stripe[456] = 24'hffffff;
assign target_only_stripe[457] = 24'hffffff;
assign target_only_stripe[458] = 24'hffffff;
assign target_only_stripe[459] = 24'hffffff;
assign target_only_stripe[460] = 24'hffffff;
assign target_only_stripe[461] = 24'hffffff;
assign target_only_stripe[462] = 24'hffffff;
assign target_only_stripe[463] = 24'h111111;
assign target_only_stripe[464] = 24'h000000;
assign target_only_stripe[465] = 24'h000000;
assign target_only_stripe[466] = 24'h000000;
assign target_only_stripe[467] = 24'h000000;
assign target_only_stripe[468] = 24'h000000;
assign target_only_stripe[469] = 24'h000000;
assign target_only_stripe[470] = 24'h000000;
assign target_only_stripe[471] = 24'h000000;
assign target_only_stripe[472] = 24'h000000;
assign target_only_stripe[473] = 24'h000000;
assign target_only_stripe[474] = 24'h000000;
assign target_only_stripe[475] = 24'h000000;
assign target_only_stripe[476] = 24'h000000;
assign target_only_stripe[477] = 24'h000000;
assign target_only_stripe[478] = 24'h000000;
assign target_only_stripe[479] = 24'h000000;
assign target_only_stripe[480] = 24'h000000;
assign target_only_stripe[481] = 24'h000000;
assign target_only_stripe[482] = 24'h000000;
assign target_only_stripe[483] = 24'h000000;
assign target_only_stripe[484] = 24'h000000;
assign target_only_stripe[485] = 24'h000000;
assign target_only_stripe[486] = 24'h000000;
assign target_only_stripe[487] = 24'h000000;
assign target_only_stripe[488] = 24'h000000;
assign target_only_stripe[489] = 24'h000000;
assign target_only_stripe[490] = 24'h000000;
assign target_only_stripe[491] = 24'h000000;
assign target_only_stripe[492] = 24'h000000;
assign target_only_stripe[493] = 24'h000000;
assign target_only_stripe[494] = 24'h000000;
assign target_only_stripe[495] = 24'h000000;
assign target_only_stripe[496] = 24'h000000;
assign target_only_stripe[497] = 24'h000000;
assign target_only_stripe[498] = 24'h000000;
assign target_only_stripe[499] = 24'h000000;
assign target_only_stripe[500] = 24'h000000;
assign target_only_stripe[501] = 24'h000000;
assign target_only_stripe[502] = 24'h000000;
assign target_only_stripe[503] = 24'h000000;
assign target_only_stripe[504] = 24'h000000;
assign target_only_stripe[505] = 24'h000000;
assign target_only_stripe[506] = 24'h000000;
assign target_only_stripe[507] = 24'h000000;
assign target_only_stripe[508] = 24'h000000;
assign target_only_stripe[509] = 24'h000000;
assign target_only_stripe[510] = 24'h000000;
assign target_only_stripe[511] = 24'h000000;
assign target_only_stripe[512] = 24'h000000;
assign target_only_stripe[513] = 24'h000000;
assign target_only_stripe[514] = 24'h000000;
assign target_only_stripe[515] = 24'h000000;
assign target_only_stripe[516] = 24'h000000;
assign target_only_stripe[517] = 24'h000000;
assign target_only_stripe[518] = 24'h000000;
assign target_only_stripe[519] = 24'h000000;
assign target_only_stripe[520] = 24'h000000;
assign target_only_stripe[521] = 24'h000000;
assign target_only_stripe[522] = 24'h000000;
assign target_only_stripe[523] = 24'h0d0d0d;
assign target_only_stripe[524] = 24'hffffff;
assign target_only_stripe[525] = 24'hffffff;
assign target_only_stripe[526] = 24'hffffff;
assign target_only_stripe[527] = 24'hffffff;
assign target_only_stripe[528] = 24'hffffff;
assign target_only_stripe[529] = 24'hffffff;
assign target_only_stripe[530] = 24'hffffff;
assign target_only_stripe[531] = 24'hffffff;
assign target_only_stripe[532] = 24'hffffff;
assign target_only_stripe[533] = 24'hffffff;
assign target_only_stripe[534] = 24'hffffff;
assign target_only_stripe[535] = 24'hffffff;
assign target_only_stripe[536] = 24'hffffff;
assign target_only_stripe[537] = 24'hffffff;
assign target_only_stripe[538] = 24'hffffff;
assign target_only_stripe[539] = 24'hffffff;
assign target_only_stripe[540] = 24'hffffff;
assign target_only_stripe[541] = 24'hffffff;
assign target_only_stripe[542] = 24'hffffff;
assign target_only_stripe[543] = 24'hffffff;
assign target_only_stripe[544] = 24'hffffff;
assign target_only_stripe[545] = 24'hffffff;
assign target_only_stripe[546] = 24'hffffff;
assign target_only_stripe[547] = 24'hffffff;
assign target_only_stripe[548] = 24'hffffff;
assign target_only_stripe[549] = 24'hffffff;
assign target_only_stripe[550] = 24'hffffff;
assign target_only_stripe[551] = 24'hffffff;
assign target_only_stripe[552] = 24'hffffff;
assign target_only_stripe[553] = 24'hffffff;
assign target_only_stripe[554] = 24'hffffff;
assign target_only_stripe[555] = 24'hffffff;
assign target_only_stripe[556] = 24'hffffff;
assign target_only_stripe[557] = 24'hffffff;
assign target_only_stripe[558] = 24'hffffff;
assign target_only_stripe[559] = 24'h010101;
assign target_only_stripe[560] = 24'h000000;
assign target_only_stripe[561] = 24'h000000;
assign target_only_stripe[562] = 24'h000000;
assign target_only_stripe[563] = 24'h000000;
assign target_only_stripe[564] = 24'h000000;
assign target_only_stripe[565] = 24'h000000;
assign target_only_stripe[566] = 24'h000000;
assign target_only_stripe[567] = 24'h000000;
assign target_only_stripe[568] = 24'h000000;
assign target_only_stripe[569] = 24'h000000;
assign target_only_stripe[570] = 24'h000000;
assign target_only_stripe[571] = 24'h000000;
assign target_only_stripe[572] = 24'h000000;
assign target_only_stripe[573] = 24'h000000;
assign target_only_stripe[574] = 24'h000000;
assign target_only_stripe[575] = 24'h000000;
assign target_only_stripe[576] = 24'h000000;
assign target_only_stripe[577] = 24'h000000;
assign target_only_stripe[578] = 24'h000000;
assign target_only_stripe[579] = 24'h000000;
assign target_only_stripe[580] = 24'h000000;
assign target_only_stripe[581] = 24'h000000;
assign target_only_stripe[582] = 24'h000000;
assign target_only_stripe[583] = 24'h000000;
assign target_only_stripe[584] = 24'h000000;
assign target_only_stripe[585] = 24'h000000;
assign target_only_stripe[586] = 24'h000000;
assign target_only_stripe[587] = 24'h000000;
assign target_only_stripe[588] = 24'h000000;
assign target_only_stripe[589] = 24'h000000;
assign target_only_stripe[590] = 24'h000000;
assign target_only_stripe[591] = 24'hcacaca;
assign target_only_stripe[592] = 24'hffffff;
assign target_only_stripe[593] = 24'hffffff;
assign target_only_stripe[594] = 24'heee4d6;
assign target_only_stripe[595] = 24'hffffff;
assign target_only_stripe[596] = 24'hffffff;
assign target_only_stripe[597] = 24'hffffff;
assign target_only_stripe[598] = 24'hffffff;
assign target_only_stripe[599] = 24'hffffff;
assign target_only_stripe[600] = 24'hffffff;
assign target_only_stripe[601] = 24'hffffff;
assign target_only_stripe[602] = 24'hffffff;
assign target_only_stripe[603] = 24'hffffff;
assign target_only_stripe[604] = 24'hffffff;
assign target_only_stripe[605] = 24'hffffff;
assign target_only_stripe[606] = 24'hffffff;
assign target_only_stripe[607] = 24'hffffff;
assign target_only_stripe[608] = 24'hffffff;
assign target_only_stripe[609] = 24'hffffff;
assign target_only_stripe[610] = 24'hffffff;
assign target_only_stripe[611] = 24'hffffff;
assign target_only_stripe[612] = 24'hffffff;
assign target_only_stripe[613] = 24'hffffff;
assign target_only_stripe[614] = 24'hffffff;
assign target_only_stripe[615] = 24'hffffff;
assign target_only_stripe[616] = 24'hffffff;
assign target_only_stripe[617] = 24'hffffff;
assign target_only_stripe[618] = 24'hffffff;
assign target_only_stripe[619] = 24'hffffff;
assign target_only_stripe[620] = 24'hffffff;
assign target_only_stripe[621] = 24'hffffff;
assign target_only_stripe[622] = 24'hffffff;
assign target_only_stripe[623] = 24'hffffff;
assign target_only_stripe[624] = 24'hffffff;
assign target_only_stripe[625] = 24'hb8b8b8;
assign target_only_stripe[626] = 24'h000000;
assign target_only_stripe[627] = 24'h000000;
assign target_only_stripe[628] = 24'h000000;
assign target_only_stripe[629] = 24'h000000;
assign target_only_stripe[630] = 24'h000000;
assign target_only_stripe[631] = 24'h000000;
assign target_only_stripe[632] = 24'h000000;
assign target_only_stripe[633] = 24'h000000;
assign target_only_stripe[634] = 24'h000000;
assign target_only_stripe[635] = 24'h000000;
assign target_only_stripe[636] = 24'h000000;
assign target_only_stripe[637] = 24'h000000;
assign target_only_stripe[638] = 24'h000000;
assign target_only_stripe[639] = 24'h000000;
assign target_only_stripe[640] = 24'h000000;
assign target_only_stripe[641] = 24'h000000;
assign target_only_stripe[642] = 24'h000000;
assign target_only_stripe[643] = 24'h000000;
assign target_only_stripe[644] = 24'h000000;
assign target_only_stripe[645] = 24'h000000;
assign target_only_stripe[646] = 24'h000000;
assign target_only_stripe[647] = 24'h000000;
assign target_only_stripe[648] = 24'h000000;
assign target_only_stripe[649] = 24'h000000;
assign target_only_stripe[650] = 24'h000000;
assign target_only_stripe[651] = 24'h000000;
assign target_only_stripe[652] = 24'h000000;
assign target_only_stripe[653] = 24'h000000;
assign target_only_stripe[654] = 24'h000000;
assign target_only_stripe[655] = 24'h000000;
assign target_only_stripe[656] = 24'h000000;
assign target_only_stripe[657] = 24'h000000;
assign target_only_stripe[658] = 24'h000000;
assign target_only_stripe[659] = 24'h000000;
assign target_only_stripe[660] = 24'h000000;
assign target_only_stripe[661] = 24'h000000;
assign target_only_stripe[662] = 24'h000000;
assign target_only_stripe[663] = 24'h000000;
assign target_only_stripe[664] = 24'h000000;
assign target_only_stripe[665] = 24'h000000;
assign target_only_stripe[666] = 24'h000000;
assign target_only_stripe[667] = 24'h000000;
assign target_only_stripe[668] = 24'h000000;
assign target_only_stripe[669] = 24'h000000;
assign target_only_stripe[670] = 24'h000000;
assign target_only_stripe[671] = 24'h000000;
assign target_only_stripe[672] = 24'h000000;
assign target_only_stripe[673] = 24'h000000;
assign target_only_stripe[674] = 24'h000000;
assign target_only_stripe[675] = 24'h000000;
assign target_only_stripe[676] = 24'h000000;
assign target_only_stripe[677] = 24'h000000;
assign target_only_stripe[678] = 24'h000000;
assign target_only_stripe[679] = 24'h000000;
assign target_only_stripe[680] = 24'h000000;
assign target_only_stripe[681] = 24'h000000;
assign target_only_stripe[682] = 24'h000000;
assign target_only_stripe[683] = 24'h000000;
assign target_only_stripe[684] = 24'h000000;
assign target_only_stripe[685] = 24'h000000;
assign target_only_stripe[686] = 24'h000000;
assign target_only_stripe[687] = 24'h000000;
assign target_only_stripe[688] = 24'h000000;
assign target_only_stripe[689] = 24'h000000;
assign target_only_stripe[690] = 24'hb9b9b9;
assign target_only_stripe[691] = 24'hffffff;
assign target_only_stripe[692] = 24'hffffff;
assign target_only_stripe[693] = 24'hffffff;
assign target_only_stripe[694] = 24'hffffff;
assign target_only_stripe[695] = 24'hffffff;
assign target_only_stripe[696] = 24'hffffff;
assign target_only_stripe[697] = 24'hffffff;
assign target_only_stripe[698] = 24'hffffff;
assign target_only_stripe[699] = 24'hffffff;
assign target_only_stripe[700] = 24'hffffff;
assign target_only_stripe[701] = 24'hffffff;
assign target_only_stripe[702] = 24'hffffff;
assign target_only_stripe[703] = 24'hffffff;
assign target_only_stripe[704] = 24'hffffff;
assign target_only_stripe[705] = 24'hffffff;
assign target_only_stripe[706] = 24'hffffff;
assign target_only_stripe[707] = 24'hffffff;
assign target_only_stripe[708] = 24'hffffff;
assign target_only_stripe[709] = 24'hffffff;
assign target_only_stripe[710] = 24'hffffff;
assign target_only_stripe[711] = 24'hffffff;
assign target_only_stripe[712] = 24'hffffff;
assign target_only_stripe[713] = 24'hfaf7f5;
assign target_only_stripe[714] = 24'hf0e8de;
assign target_only_stripe[715] = 24'hffffff;
assign target_only_stripe[716] = 24'hffffff;
assign target_only_stripe[717] = 24'hffffff;
assign target_only_stripe[718] = 24'hffffff;
assign target_only_stripe[719] = 24'hffffff;
assign target_only_stripe[720] = 24'hffffff;
assign target_only_stripe[721] = 24'hffffff;
assign target_only_stripe[722] = 24'hffffff;
assign target_only_stripe[723] = 24'he6e1df;
assign target_only_stripe[724] = 24'h262626;
assign target_only_stripe[725] = 24'h000000;
assign target_only_stripe[726] = 24'h000000;
assign target_only_stripe[727] = 24'h000000;
assign target_only_stripe[728] = 24'h000000;
assign target_only_stripe[729] = 24'h000000;
assign target_only_stripe[730] = 24'h000000;
assign target_only_stripe[731] = 24'h000000;
assign target_only_stripe[732] = 24'h000000;
assign target_only_stripe[733] = 24'h000000;
assign target_only_stripe[734] = 24'h000000;
assign target_only_stripe[735] = 24'h000000;
assign target_only_stripe[736] = 24'h000000;
assign target_only_stripe[737] = 24'h000000;
assign target_only_stripe[738] = 24'h000000;
assign target_only_stripe[739] = 24'h000000;
assign target_only_stripe[740] = 24'h000000;
assign target_only_stripe[741] = 24'h000000;
assign target_only_stripe[742] = 24'h000000;
assign target_only_stripe[743] = 24'h000000;
assign target_only_stripe[744] = 24'h000000;
assign target_only_stripe[745] = 24'h000000;
assign target_only_stripe[746] = 24'h000000;
assign target_only_stripe[747] = 24'h000000;
assign target_only_stripe[748] = 24'h000000;
assign target_only_stripe[749] = 24'h000000;
assign target_only_stripe[750] = 24'h000000;
assign target_only_stripe[751] = 24'h000000;
assign target_only_stripe[752] = 24'h000000;
assign target_only_stripe[753] = 24'h000000;
assign target_only_stripe[754] = 24'h000000;
assign target_only_stripe[755] = 24'h000000;
assign target_only_stripe[756] = 24'h1c1c1c;
assign target_only_stripe[757] = 24'hffffff;
assign target_only_stripe[758] = 24'hffffff;
assign target_only_stripe[759] = 24'hffffff;
assign target_only_stripe[760] = 24'hffffff;
assign target_only_stripe[761] = 24'hffffff;
assign target_only_stripe[762] = 24'hffffff;
assign target_only_stripe[763] = 24'hffffff;
assign target_only_stripe[764] = 24'hffffff;
assign target_only_stripe[765] = 24'hffffff;
assign target_only_stripe[766] = 24'hffffff;
assign target_only_stripe[767] = 24'hffffff;
assign target_only_stripe[768] = 24'hffffff;
assign target_only_stripe[769] = 24'hffffff;
assign target_only_stripe[770] = 24'hffffff;
assign target_only_stripe[771] = 24'hffffff;
assign target_only_stripe[772] = 24'hffffff;
assign target_only_stripe[773] = 24'hffffff;
assign target_only_stripe[774] = 24'hffffff;
assign target_only_stripe[775] = 24'hffffff;
assign target_only_stripe[776] = 24'hffffff;
assign target_only_stripe[777] = 24'hffffff;
assign target_only_stripe[778] = 24'hffffff;
assign target_only_stripe[779] = 24'hffffff;
assign target_only_stripe[780] = 24'hffffff;
assign target_only_stripe[781] = 24'hffffff;
assign target_only_stripe[782] = 24'hffffff;
assign target_only_stripe[783] = 24'hffffff;
assign target_only_stripe[784] = 24'hffffff;
assign target_only_stripe[785] = 24'hffffff;
assign target_only_stripe[786] = 24'hffffff;
assign target_only_stripe[787] = 24'hffffff;
assign target_only_stripe[788] = 24'hffffff;
assign target_only_stripe[789] = 24'hffffff;
assign target_only_stripe[790] = 24'hffffff;
assign target_only_stripe[791] = 24'h9d9d9d;
assign target_only_stripe[792] = 24'h000000;
assign target_only_stripe[793] = 24'h000000;
assign target_only_stripe[794] = 24'h000000;
assign target_only_stripe[795] = 24'h000000;
assign target_only_stripe[796] = 24'h000000;
assign target_only_stripe[797] = 24'h000000;
assign target_only_stripe[798] = 24'h000000;
assign target_only_stripe[799] = 24'h000000;
assign target_only_stripe[800] = 24'h000000;
assign target_only_stripe[801] = 24'h000000;
assign target_only_stripe[802] = 24'h000000;
assign target_only_stripe[803] = 24'h000000;
assign target_only_stripe[804] = 24'h000000;
assign target_only_stripe[805] = 24'h000000;
assign target_only_stripe[806] = 24'h000000;
assign target_only_stripe[807] = 24'h000000;
assign target_only_stripe[808] = 24'h000000;
assign target_only_stripe[809] = 24'h000000;
assign target_only_stripe[810] = 24'h000000;
assign target_only_stripe[811] = 24'h000000;
assign target_only_stripe[812] = 24'h000000;
assign target_only_stripe[813] = 24'h000000;
assign target_only_stripe[814] = 24'h000000;
assign target_only_stripe[815] = 24'h000000;
assign target_only_stripe[816] = 24'h000000;
assign target_only_stripe[817] = 24'h000000;
assign target_only_stripe[818] = 24'h000000;
assign target_only_stripe[819] = 24'h000000;
assign target_only_stripe[820] = 24'h000000;
assign target_only_stripe[821] = 24'h000000;
assign target_only_stripe[822] = 24'h000000;
assign target_only_stripe[823] = 24'h000000;
assign target_only_stripe[824] = 24'h000000;
assign target_only_stripe[825] = 24'h000000;
assign target_only_stripe[826] = 24'h000000;
assign target_only_stripe[827] = 24'h000000;
assign target_only_stripe[828] = 24'h000000;
assign target_only_stripe[829] = 24'h000000;
assign target_only_stripe[830] = 24'h000000;
assign target_only_stripe[831] = 24'h000000;
assign target_only_stripe[832] = 24'h000000;
assign target_only_stripe[833] = 24'h000000;
assign target_only_stripe[834] = 24'h000000;
assign target_only_stripe[835] = 24'h000000;
assign target_only_stripe[836] = 24'h000000;
assign target_only_stripe[837] = 24'h000000;
assign target_only_stripe[838] = 24'h000000;
assign target_only_stripe[839] = 24'h000000;
assign target_only_stripe[840] = 24'h000000;
assign target_only_stripe[841] = 24'h000000;
assign target_only_stripe[842] = 24'h000000;
assign target_only_stripe[843] = 24'h000000;
assign target_only_stripe[844] = 24'h000000;
assign target_only_stripe[845] = 24'h000000;
assign target_only_stripe[846] = 24'h000000;
assign target_only_stripe[847] = 24'h000000;
assign target_only_stripe[848] = 24'h000000;
assign target_only_stripe[849] = 24'h000000;
assign target_only_stripe[850] = 24'h000000;
assign target_only_stripe[851] = 24'h000000;
assign target_only_stripe[852] = 24'h000000;
assign target_only_stripe[853] = 24'h969696;
assign target_only_stripe[854] = 24'hffffff;
assign target_only_stripe[855] = 24'hffffff;
assign target_only_stripe[856] = 24'hffffff;
assign target_only_stripe[857] = 24'hffffff;
assign target_only_stripe[858] = 24'hffffff;
assign target_only_stripe[859] = 24'hffffff;
assign target_only_stripe[860] = 24'hffffff;
assign target_only_stripe[861] = 24'hffffff;
assign target_only_stripe[862] = 24'hffffff;
assign target_only_stripe[863] = 24'hffffff;
assign target_only_stripe[864] = 24'hffffff;
assign target_only_stripe[865] = 24'hffffff;
assign target_only_stripe[866] = 24'hffffff;
assign target_only_stripe[867] = 24'hffffff;
assign target_only_stripe[868] = 24'hffffff;
assign target_only_stripe[869] = 24'hffffff;
assign target_only_stripe[870] = 24'hffffff;
assign target_only_stripe[871] = 24'hffffff;
assign target_only_stripe[872] = 24'hffffff;
assign target_only_stripe[873] = 24'hffffff;
assign target_only_stripe[874] = 24'hffffff;
assign target_only_stripe[875] = 24'hffffff;
assign target_only_stripe[876] = 24'hffffff;
assign target_only_stripe[877] = 24'hffffff;
assign target_only_stripe[878] = 24'hffffff;
assign target_only_stripe[879] = 24'hffffff;
assign target_only_stripe[880] = 24'hffffff;
assign target_only_stripe[881] = 24'hffffff;
assign target_only_stripe[882] = 24'hffffff;
assign target_only_stripe[883] = 24'hffffff;
assign target_only_stripe[884] = 24'hffffff;
assign target_only_stripe[885] = 24'hffffff;
assign target_only_stripe[886] = 24'hffffff;
assign target_only_stripe[887] = 24'hffffff;
assign target_only_stripe[888] = 24'h222222;
assign target_only_stripe[889] = 24'h000000;
assign target_only_stripe[890] = 24'h000000;
assign target_only_stripe[891] = 24'h000000;
assign target_only_stripe[892] = 24'h000000;
assign target_only_stripe[893] = 24'h000000;
assign target_only_stripe[894] = 24'h000000;
assign target_only_stripe[895] = 24'h000000;
assign target_only_stripe[896] = 24'h000000;
assign target_only_stripe[897] = 24'h000000;
assign target_only_stripe[898] = 24'h000000;
assign target_only_stripe[899] = 24'h000000;
assign target_only_stripe[900] = 24'h000000;
assign target_only_stripe[901] = 24'h000000;
assign target_only_stripe[902] = 24'h000000;
assign target_only_stripe[903] = 24'h000000;
assign target_only_stripe[904] = 24'h000000;
assign target_only_stripe[905] = 24'h000000;
assign target_only_stripe[906] = 24'h000000;
assign target_only_stripe[907] = 24'h000000;
assign target_only_stripe[908] = 24'h000000;
assign target_only_stripe[909] = 24'h000000;
assign target_only_stripe[910] = 24'h000000;
assign target_only_stripe[911] = 24'h000000;
assign target_only_stripe[912] = 24'h000000;
assign target_only_stripe[913] = 24'h000000;
assign target_only_stripe[914] = 24'h000000;
assign target_only_stripe[915] = 24'h000000;
assign target_only_stripe[916] = 24'h000000;
assign target_only_stripe[917] = 24'h000000;
assign target_only_stripe[918] = 24'h000000;
assign target_only_stripe[919] = 24'h000000;
assign target_only_stripe[920] = 24'h1d1d1d;
assign target_only_stripe[921] = 24'he7e7e7;
assign target_only_stripe[922] = 24'hffffff;
assign target_only_stripe[923] = 24'hf0e8de;
assign target_only_stripe[924] = 24'hfaf7f5;
assign target_only_stripe[925] = 24'hffffff;
assign target_only_stripe[926] = 24'hffffff;
assign target_only_stripe[927] = 24'hffffff;
assign target_only_stripe[928] = 24'hffffff;
assign target_only_stripe[929] = 24'hffffff;
assign target_only_stripe[930] = 24'hffffff;
assign target_only_stripe[931] = 24'hffffff;
assign target_only_stripe[932] = 24'hffffff;
assign target_only_stripe[933] = 24'hffffff;
assign target_only_stripe[934] = 24'hffffff;
assign target_only_stripe[935] = 24'hffffff;
assign target_only_stripe[936] = 24'hffffff;
assign target_only_stripe[937] = 24'hffffff;
assign target_only_stripe[938] = 24'hffffff;
assign target_only_stripe[939] = 24'hffffff;
assign target_only_stripe[940] = 24'hffffff;
assign target_only_stripe[941] = 24'hffffff;
assign target_only_stripe[942] = 24'hffffff;
assign target_only_stripe[943] = 24'hffffff;
assign target_only_stripe[944] = 24'hffffff;
assign target_only_stripe[945] = 24'hffffff;
assign target_only_stripe[946] = 24'hffffff;
assign target_only_stripe[947] = 24'hffffff;
assign target_only_stripe[948] = 24'hffffff;
assign target_only_stripe[949] = 24'hffffff;
assign target_only_stripe[950] = 24'hffffff;
assign target_only_stripe[951] = 24'hffffff;
assign target_only_stripe[952] = 24'hffffff;
assign target_only_stripe[953] = 24'hffffff;
assign target_only_stripe[954] = 24'hbfbfbf;
assign target_only_stripe[955] = 24'h000000;
assign target_only_stripe[956] = 24'h000000;
assign target_only_stripe[957] = 24'h000000;
assign target_only_stripe[958] = 24'h000000;
assign target_only_stripe[959] = 24'h000000;
assign target_only_stripe[960] = 24'h000000;
assign target_only_stripe[961] = 24'h000000;
assign target_only_stripe[962] = 24'h000000;
assign target_only_stripe[963] = 24'h000000;
assign target_only_stripe[964] = 24'h000000;
assign target_only_stripe[965] = 24'h000000;
assign target_only_stripe[966] = 24'h000000;
assign target_only_stripe[967] = 24'h000000;
assign target_only_stripe[968] = 24'h000000;
assign target_only_stripe[969] = 24'h000000;
assign target_only_stripe[970] = 24'h000000;
assign target_only_stripe[971] = 24'h000000;
assign target_only_stripe[972] = 24'h000000;
assign target_only_stripe[973] = 24'h000000;
assign target_only_stripe[974] = 24'h000000;
assign target_only_stripe[975] = 24'h000000;
assign target_only_stripe[976] = 24'h000000;
assign target_only_stripe[977] = 24'h000000;
assign target_only_stripe[978] = 24'h000000;
assign target_only_stripe[979] = 24'h000000;
assign target_only_stripe[980] = 24'h000000;
assign target_only_stripe[981] = 24'h000000;
assign target_only_stripe[982] = 24'h000000;
assign target_only_stripe[983] = 24'h000000;
assign target_only_stripe[984] = 24'h000000;
assign target_only_stripe[985] = 24'h000000;
assign target_only_stripe[986] = 24'h000000;
assign target_only_stripe[987] = 24'h000000;
assign target_only_stripe[988] = 24'h000000;
assign target_only_stripe[989] = 24'h000000;
assign target_only_stripe[990] = 24'h000000;
assign target_only_stripe[991] = 24'h000000;
assign target_only_stripe[992] = 24'h000000;
assign target_only_stripe[993] = 24'h000000;
assign target_only_stripe[994] = 24'h000000;
assign target_only_stripe[995] = 24'h000000;
assign target_only_stripe[996] = 24'h000000;
assign target_only_stripe[997] = 24'h000000;
assign target_only_stripe[998] = 24'h000000;
assign target_only_stripe[999] = 24'h000000;
assign target_only_stripe[1000] = 24'h000000;
assign target_only_stripe[1001] = 24'h000000;
assign target_only_stripe[1002] = 24'h000000;
assign target_only_stripe[1003] = 24'h000000;
assign target_only_stripe[1004] = 24'h000000;
assign target_only_stripe[1005] = 24'h000000;
assign target_only_stripe[1006] = 24'h000000;
assign target_only_stripe[1007] = 24'h000000;
assign target_only_stripe[1008] = 24'h000000;
assign target_only_stripe[1009] = 24'h000000;
assign target_only_stripe[1010] = 24'h000000;
assign target_only_stripe[1011] = 24'h000000;
assign target_only_stripe[1012] = 24'h000000;
assign target_only_stripe[1013] = 24'h000000;
assign target_only_stripe[1014] = 24'h000000;
assign target_only_stripe[1015] = 24'h000000;
assign target_only_stripe[1016] = 24'h000000;
assign target_only_stripe[1017] = 24'h000000;
assign target_only_stripe[1018] = 24'h010101;
assign target_only_stripe[1019] = 24'hbdbdbd;
assign target_only_stripe[1020] = 24'hffffff;
assign target_only_stripe[1021] = 24'hffffff;
assign target_only_stripe[1022] = 24'hffffff;
assign target_only_stripe[1023] = 24'hffffff;
assign target_only_stripe[1024] = 24'hffffff;
assign target_only_stripe[1025] = 24'hffffff;
assign target_only_stripe[1026] = 24'hffffff;
assign target_only_stripe[1027] = 24'hffffff;
assign target_only_stripe[1028] = 24'hffffff;
assign target_only_stripe[1029] = 24'hffffff;
assign target_only_stripe[1030] = 24'hffffff;
assign target_only_stripe[1031] = 24'hffffff;
assign target_only_stripe[1032] = 24'hffffff;
assign target_only_stripe[1033] = 24'hffffff;
assign target_only_stripe[1034] = 24'hffffff;
assign target_only_stripe[1035] = 24'hffffff;
assign target_only_stripe[1036] = 24'hffffff;
assign target_only_stripe[1037] = 24'hffffff;
assign target_only_stripe[1038] = 24'hffffff;
assign target_only_stripe[1039] = 24'hffffff;
assign target_only_stripe[1040] = 24'hffffff;
assign target_only_stripe[1041] = 24'hffffff;
assign target_only_stripe[1042] = 24'hffffff;
assign target_only_stripe[1043] = 24'hffffff;
assign target_only_stripe[1044] = 24'hffffff;
assign target_only_stripe[1045] = 24'hffffff;
assign target_only_stripe[1046] = 24'hffffff;
assign target_only_stripe[1047] = 24'hffffff;
assign target_only_stripe[1048] = 24'hffffff;
assign target_only_stripe[1049] = 24'hffffff;
assign target_only_stripe[1050] = 24'hffffff;
assign target_only_stripe[1051] = 24'hffffff;
assign target_only_stripe[1052] = 24'hdedede;
assign target_only_stripe[1053] = 24'h1b1b1b;
assign target_only_stripe[1054] = 24'h000000;
assign target_only_stripe[1055] = 24'h000000;
assign target_only_stripe[1056] = 24'h000000;
assign target_only_stripe[1057] = 24'h000000;
assign target_only_stripe[1058] = 24'h000000;
assign target_only_stripe[1059] = 24'h000000;
assign target_only_stripe[1060] = 24'h000000;
assign target_only_stripe[1061] = 24'h000000;
assign target_only_stripe[1062] = 24'h000000;
assign target_only_stripe[1063] = 24'h000000;
assign target_only_stripe[1064] = 24'h000000;
assign target_only_stripe[1065] = 24'h000000;
assign target_only_stripe[1066] = 24'h000000;
assign target_only_stripe[1067] = 24'h000000;
assign target_only_stripe[1068] = 24'h000000;
assign target_only_stripe[1069] = 24'h000000;
assign target_only_stripe[1070] = 24'h000000;
assign target_only_stripe[1071] = 24'h000000;
assign target_only_stripe[1072] = 24'h000000;
assign target_only_stripe[1073] = 24'h000000;
assign target_only_stripe[1074] = 24'h000000;
assign target_only_stripe[1075] = 24'h000000;
assign target_only_stripe[1076] = 24'h000000;
assign target_only_stripe[1077] = 24'h000000;
assign target_only_stripe[1078] = 24'h000000;
assign target_only_stripe[1079] = 24'h000000;
assign target_only_stripe[1080] = 24'h000000;
assign target_only_stripe[1081] = 24'h000000;
assign target_only_stripe[1082] = 24'h000000;
assign target_only_stripe[1083] = 24'h000000;
assign target_only_stripe[1084] = 24'h000000;
assign target_only_stripe[1085] = 24'h2f2f2f;
assign target_only_stripe[1086] = 24'hffffff;
assign target_only_stripe[1087] = 24'hffffff;
assign target_only_stripe[1088] = 24'hffffff;
assign target_only_stripe[1089] = 24'hffffff;
assign target_only_stripe[1090] = 24'hffffff;
assign target_only_stripe[1091] = 24'hffffff;
assign target_only_stripe[1092] = 24'hffffff;
assign target_only_stripe[1093] = 24'hffffff;
assign target_only_stripe[1094] = 24'hffffff;
assign target_only_stripe[1095] = 24'hffffff;
assign target_only_stripe[1096] = 24'hffffff;
assign target_only_stripe[1097] = 24'hffffff;
assign target_only_stripe[1098] = 24'hffffff;
assign target_only_stripe[1099] = 24'hffffff;
assign target_only_stripe[1100] = 24'hffffff;
assign target_only_stripe[1101] = 24'hffffff;
assign target_only_stripe[1102] = 24'hffffff;
assign target_only_stripe[1103] = 24'hffffff;
assign target_only_stripe[1104] = 24'hffffff;
assign target_only_stripe[1105] = 24'hffffff;
assign target_only_stripe[1106] = 24'hffffff;
assign target_only_stripe[1107] = 24'hffffff;
assign target_only_stripe[1108] = 24'hffffff;
assign target_only_stripe[1109] = 24'hffffff;
assign target_only_stripe[1110] = 24'hffffff;
assign target_only_stripe[1111] = 24'hffffff;
assign target_only_stripe[1112] = 24'hffffff;
assign target_only_stripe[1113] = 24'hffffff;
assign target_only_stripe[1114] = 24'hffffff;
assign target_only_stripe[1115] = 24'hffffff;
assign target_only_stripe[1116] = 24'hffffff;
assign target_only_stripe[1117] = 24'hffffff;
assign target_only_stripe[1118] = 24'hffffff;
assign target_only_stripe[1119] = 24'hffffff;
assign target_only_stripe[1120] = 24'hffffff;
assign target_only_stripe[1121] = 24'h000000;
assign target_only_stripe[1122] = 24'h000000;
assign target_only_stripe[1123] = 24'h000000;
assign target_only_stripe[1124] = 24'h000000;
assign target_only_stripe[1125] = 24'h000000;
assign target_only_stripe[1126] = 24'h000000;
assign target_only_stripe[1127] = 24'h000000;
assign target_only_stripe[1128] = 24'h000000;
assign target_only_stripe[1129] = 24'h000000;
assign target_only_stripe[1130] = 24'h000000;
assign target_only_stripe[1131] = 24'h000000;
assign target_only_stripe[1132] = 24'h000000;
assign target_only_stripe[1133] = 24'h000000;
assign target_only_stripe[1134] = 24'h000000;
assign target_only_stripe[1135] = 24'h000000;
assign target_only_stripe[1136] = 24'h000000;
assign target_only_stripe[1137] = 24'h000000;
assign target_only_stripe[1138] = 24'h000000;
assign target_only_stripe[1139] = 24'h000000;
assign target_only_stripe[1140] = 24'h000000;
assign target_only_stripe[1141] = 24'h000000;
assign target_only_stripe[1142] = 24'h000000;
assign target_only_stripe[1143] = 24'h000000;
assign target_only_stripe[1144] = 24'h000000;
assign target_only_stripe[1145] = 24'h000000;
assign target_only_stripe[1146] = 24'h000000;
assign target_only_stripe[1147] = 24'h000000;
assign target_only_stripe[1148] = 24'h000000;
assign target_only_stripe[1149] = 24'h000000;
assign target_only_stripe[1150] = 24'h000000;
assign target_only_stripe[1151] = 24'h000000;
assign target_only_stripe[1152] = 24'h000000;
assign target_only_stripe[1153] = 24'h000000;
assign target_only_stripe[1154] = 24'h000000;
assign target_only_stripe[1155] = 24'h000000;
assign target_only_stripe[1156] = 24'h000000;
assign target_only_stripe[1157] = 24'h000000;
assign target_only_stripe[1158] = 24'h000000;
assign target_only_stripe[1159] = 24'h000000;
assign target_only_stripe[1160] = 24'h000000;
assign target_only_stripe[1161] = 24'h000000;
assign target_only_stripe[1162] = 24'h000000;
assign target_only_stripe[1163] = 24'h000000;
assign target_only_stripe[1164] = 24'h000000;
assign target_only_stripe[1165] = 24'h000000;
assign target_only_stripe[1166] = 24'h000000;
assign target_only_stripe[1167] = 24'h000000;
assign target_only_stripe[1168] = 24'h000000;
assign target_only_stripe[1169] = 24'h000000;
assign target_only_stripe[1170] = 24'h000000;
assign target_only_stripe[1171] = 24'h000000;
assign target_only_stripe[1172] = 24'h000000;
assign target_only_stripe[1173] = 24'h000000;
assign target_only_stripe[1174] = 24'h000000;
assign target_only_stripe[1175] = 24'h000000;
assign target_only_stripe[1176] = 24'h000000;
assign target_only_stripe[1177] = 24'h000000;
assign target_only_stripe[1178] = 24'h000000;
assign target_only_stripe[1179] = 24'h000000;
assign target_only_stripe[1180] = 24'h000000;
assign target_only_stripe[1181] = 24'h000000;
assign target_only_stripe[1182] = 24'h818181;
assign target_only_stripe[1183] = 24'hffffff;
assign target_only_stripe[1184] = 24'hffffff;
assign target_only_stripe[1185] = 24'hffffff;
assign target_only_stripe[1186] = 24'hffffff;
assign target_only_stripe[1187] = 24'hffffff;
assign target_only_stripe[1188] = 24'hffffff;
assign target_only_stripe[1189] = 24'hffffff;
assign target_only_stripe[1190] = 24'hffffff;
assign target_only_stripe[1191] = 24'hffffff;
assign target_only_stripe[1192] = 24'hffffff;
assign target_only_stripe[1193] = 24'hffffff;
assign target_only_stripe[1194] = 24'hffffff;
assign target_only_stripe[1195] = 24'hffffff;
assign target_only_stripe[1196] = 24'hffffff;
assign target_only_stripe[1197] = 24'hffffff;
assign target_only_stripe[1198] = 24'hffffff;
assign target_only_stripe[1199] = 24'hffffff;
assign target_only_stripe[1200] = 24'hffffff;
assign target_only_stripe[1201] = 24'hffffff;
assign target_only_stripe[1202] = 24'hffffff;
assign target_only_stripe[1203] = 24'hffffff;
assign target_only_stripe[1204] = 24'hffffff;
assign target_only_stripe[1205] = 24'hffffff;
assign target_only_stripe[1206] = 24'hffffff;
assign target_only_stripe[1207] = 24'hffffff;
assign target_only_stripe[1208] = 24'hffffff;
assign target_only_stripe[1209] = 24'hffffff;
assign target_only_stripe[1210] = 24'hffffff;
assign target_only_stripe[1211] = 24'hffffff;
assign target_only_stripe[1212] = 24'hffffff;
assign target_only_stripe[1213] = 24'hffffff;
assign target_only_stripe[1214] = 24'hffffff;
assign target_only_stripe[1215] = 24'hffffff;
assign target_only_stripe[1216] = 24'hffffff;
assign target_only_stripe[1217] = 24'h383838;
assign target_only_stripe[1218] = 24'h000000;
assign target_only_stripe[1219] = 24'h000000;
assign target_only_stripe[1220] = 24'h000000;
assign target_only_stripe[1221] = 24'h000000;
assign target_only_stripe[1222] = 24'h000000;
assign target_only_stripe[1223] = 24'h000000;
assign target_only_stripe[1224] = 24'h000000;
assign target_only_stripe[1225] = 24'h000000;
assign target_only_stripe[1226] = 24'h000000;
assign target_only_stripe[1227] = 24'h000000;
assign target_only_stripe[1228] = 24'h000000;
assign target_only_stripe[1229] = 24'h000000;
assign target_only_stripe[1230] = 24'h000000;
assign target_only_stripe[1231] = 24'h000000;
assign target_only_stripe[1232] = 24'h000000;
assign target_only_stripe[1233] = 24'h000000;
assign target_only_stripe[1234] = 24'h000000;
assign target_only_stripe[1235] = 24'h000000;
assign target_only_stripe[1236] = 24'h000000;
assign target_only_stripe[1237] = 24'h000000;
assign target_only_stripe[1238] = 24'h000000;
assign target_only_stripe[1239] = 24'h000000;
assign target_only_stripe[1240] = 24'h000000;
assign target_only_stripe[1241] = 24'h000000;
assign target_only_stripe[1242] = 24'h000000;
assign target_only_stripe[1243] = 24'h000000;
assign target_only_stripe[1244] = 24'h000000;
assign target_only_stripe[1245] = 24'h000000;
assign target_only_stripe[1246] = 24'h000000;
assign target_only_stripe[1247] = 24'h000000;
assign target_only_stripe[1248] = 24'h000000;
assign target_only_stripe[1249] = 24'h131313;
assign target_only_stripe[1250] = 24'hd9d9d9;
assign target_only_stripe[1251] = 24'hffffff;
assign target_only_stripe[1252] = 24'heee4d6;
assign target_only_stripe[1253] = 24'hfaf7f5;
assign target_only_stripe[1254] = 24'hffffff;
assign target_only_stripe[1255] = 24'hffffff;
assign target_only_stripe[1256] = 24'hffffff;
assign target_only_stripe[1257] = 24'hffffff;
assign target_only_stripe[1258] = 24'hffffff;
assign target_only_stripe[1259] = 24'hffffff;
assign target_only_stripe[1260] = 24'hffffff;
assign target_only_stripe[1261] = 24'hffffff;
assign target_only_stripe[1262] = 24'hffffff;
assign target_only_stripe[1263] = 24'hffffff;
assign target_only_stripe[1264] = 24'hffffff;
assign target_only_stripe[1265] = 24'hffffff;
assign target_only_stripe[1266] = 24'hffffff;
assign target_only_stripe[1267] = 24'hffffff;
assign target_only_stripe[1268] = 24'hffffff;
assign target_only_stripe[1269] = 24'hffffff;
assign target_only_stripe[1270] = 24'hffffff;
assign target_only_stripe[1271] = 24'hffffff;
assign target_only_stripe[1272] = 24'hffffff;
assign target_only_stripe[1273] = 24'hffffff;
assign target_only_stripe[1274] = 24'hffffff;
assign target_only_stripe[1275] = 24'hffffff;
assign target_only_stripe[1276] = 24'hffffff;
assign target_only_stripe[1277] = 24'hffffff;
assign target_only_stripe[1278] = 24'hffffff;
assign target_only_stripe[1279] = 24'hffffff;
assign target_only_stripe[1280] = 24'hffffff;
assign target_only_stripe[1281] = 24'hffffff;
assign target_only_stripe[1282] = 24'hffffff;
assign target_only_stripe[1283] = 24'hc3c3c3;
assign target_only_stripe[1284] = 24'h010101;
assign target_only_stripe[1285] = 24'h000000;
assign target_only_stripe[1286] = 24'h000000;
assign target_only_stripe[1287] = 24'h000000;
assign target_only_stripe[1288] = 24'h000000;
assign target_only_stripe[1289] = 24'h000000;
assign target_only_stripe[1290] = 24'h000000;
assign target_only_stripe[1291] = 24'h000000;
assign target_only_stripe[1292] = 24'h000000;
assign target_only_stripe[1293] = 24'h000000;
assign target_only_stripe[1294] = 24'h000000;
assign target_only_stripe[1295] = 24'h000000;
assign target_only_stripe[1296] = 24'h000000;
assign target_only_stripe[1297] = 24'h000000;
assign target_only_stripe[1298] = 24'h000000;
assign target_only_stripe[1299] = 24'h000000;
assign target_only_stripe[1300] = 24'h000000;
assign target_only_stripe[1301] = 24'h000000;
assign target_only_stripe[1302] = 24'h000000;
assign target_only_stripe[1303] = 24'h000000;
assign target_only_stripe[1304] = 24'h000000;
assign target_only_stripe[1305] = 24'h000000;
assign target_only_stripe[1306] = 24'h000000;
assign target_only_stripe[1307] = 24'h000000;
assign target_only_stripe[1308] = 24'h000000;
assign target_only_stripe[1309] = 24'h000000;
assign target_only_stripe[1310] = 24'h000000;
assign target_only_stripe[1311] = 24'h000000;
assign target_only_stripe[1312] = 24'h000000;
assign target_only_stripe[1313] = 24'h000000;
assign target_only_stripe[1314] = 24'h000000;
assign target_only_stripe[1315] = 24'h000000;
assign target_only_stripe[1316] = 24'h000000;
assign target_only_stripe[1317] = 24'h000000;
assign target_only_stripe[1318] = 24'h000000;
assign target_only_stripe[1319] = 24'h000000;
assign target_only_stripe[1320] = 24'h000000;
assign target_only_stripe[1321] = 24'h000000;
assign target_only_stripe[1322] = 24'h000000;
assign target_only_stripe[1323] = 24'h000000;
assign target_only_stripe[1324] = 24'h000000;
assign target_only_stripe[1325] = 24'h000000;
assign target_only_stripe[1326] = 24'h000000;
assign target_only_stripe[1327] = 24'h000000;
assign target_only_stripe[1328] = 24'h000000;
assign target_only_stripe[1329] = 24'h000000;
assign target_only_stripe[1330] = 24'h000000;
assign target_only_stripe[1331] = 24'h000000;
assign target_only_stripe[1332] = 24'h000000;
assign target_only_stripe[1333] = 24'h000000;
assign target_only_stripe[1334] = 24'h000000;
assign target_only_stripe[1335] = 24'h000000;
assign target_only_stripe[1336] = 24'h000000;
assign target_only_stripe[1337] = 24'h000000;
assign target_only_stripe[1338] = 24'h000000;
assign target_only_stripe[1339] = 24'h000000;
assign target_only_stripe[1340] = 24'h000000;
assign target_only_stripe[1341] = 24'h000000;
assign target_only_stripe[1342] = 24'h000000;
assign target_only_stripe[1343] = 24'h000000;
assign target_only_stripe[1344] = 24'h000000;
assign target_only_stripe[1345] = 24'h000000;
assign target_only_stripe[1346] = 24'h000000;
assign target_only_stripe[1347] = 24'h070707;
assign target_only_stripe[1348] = 24'hcdcdcd;
assign target_only_stripe[1349] = 24'hffffff;
assign target_only_stripe[1350] = 24'hffffff;
assign target_only_stripe[1351] = 24'hffffff;
assign target_only_stripe[1352] = 24'hffffff;
assign target_only_stripe[1353] = 24'hffffff;
assign target_only_stripe[1354] = 24'hffffff;
assign target_only_stripe[1355] = 24'hffffff;
assign target_only_stripe[1356] = 24'hffffff;
assign target_only_stripe[1357] = 24'hffffff;
assign target_only_stripe[1358] = 24'hffffff;
assign target_only_stripe[1359] = 24'hffffff;
assign target_only_stripe[1360] = 24'hffffff;
assign target_only_stripe[1361] = 24'hffffff;
assign target_only_stripe[1362] = 24'hffffff;
assign target_only_stripe[1363] = 24'hffffff;
assign target_only_stripe[1364] = 24'hffffff;
assign target_only_stripe[1365] = 24'hffffff;
assign target_only_stripe[1366] = 24'hffffff;
assign target_only_stripe[1367] = 24'hffffff;
assign target_only_stripe[1368] = 24'hffffff;
assign target_only_stripe[1369] = 24'hffffff;
assign target_only_stripe[1370] = 24'hffffff;
assign target_only_stripe[1371] = 24'hffffff;
assign target_only_stripe[1372] = 24'hffffff;
assign target_only_stripe[1373] = 24'hffffff;
assign target_only_stripe[1374] = 24'hffffff;
assign target_only_stripe[1375] = 24'hffffff;
assign target_only_stripe[1376] = 24'hffffff;
assign target_only_stripe[1377] = 24'hffffff;
assign target_only_stripe[1378] = 24'hffffff;
assign target_only_stripe[1379] = 24'hffffff;
assign target_only_stripe[1380] = 24'hffffff;
assign target_only_stripe[1381] = 24'hd3d3d3;
assign target_only_stripe[1382] = 24'h101010;
assign target_only_stripe[1383] = 24'h000000;
assign target_only_stripe[1384] = 24'h000000;
assign target_only_stripe[1385] = 24'h000000;
assign target_only_stripe[1386] = 24'h000000;
assign target_only_stripe[1387] = 24'h000000;
assign target_only_stripe[1388] = 24'h000000;
assign target_only_stripe[1389] = 24'h000000;
assign target_only_stripe[1390] = 24'h000000;
assign target_only_stripe[1391] = 24'h000000;
assign target_only_stripe[1392] = 24'h000000;
assign target_only_stripe[1393] = 24'h000000;
assign target_only_stripe[1394] = 24'h000000;
assign target_only_stripe[1395] = 24'h000000;
assign target_only_stripe[1396] = 24'h000000;
assign target_only_stripe[1397] = 24'h000000;
assign target_only_stripe[1398] = 24'h000000;
assign target_only_stripe[1399] = 24'h000000;
assign target_only_stripe[1400] = 24'h000000;
assign target_only_stripe[1401] = 24'h000000;
assign target_only_stripe[1402] = 24'h000000;
assign target_only_stripe[1403] = 24'h000000;
assign target_only_stripe[1404] = 24'h000000;
assign target_only_stripe[1405] = 24'h000000;
assign target_only_stripe[1406] = 24'h000000;
assign target_only_stripe[1407] = 24'h000000;
assign target_only_stripe[1408] = 24'h000000;
assign target_only_stripe[1409] = 24'h000000;
assign target_only_stripe[1410] = 24'h000000;
assign target_only_stripe[1411] = 24'h000000;
assign target_only_stripe[1412] = 24'h000000;
assign target_only_stripe[1413] = 24'h000000;
assign target_only_stripe[1414] = 24'h393939;
assign target_only_stripe[1415] = 24'hffffff;
assign target_only_stripe[1416] = 24'hffffff;
assign target_only_stripe[1417] = 24'hffffff;
assign target_only_stripe[1418] = 24'hffffff;
assign target_only_stripe[1419] = 24'hffffff;
assign target_only_stripe[1420] = 24'hffffff;
assign target_only_stripe[1421] = 24'hffffff;
assign target_only_stripe[1422] = 24'hffffff;
assign target_only_stripe[1423] = 24'hffffff;
assign target_only_stripe[1424] = 24'hffffff;
assign target_only_stripe[1425] = 24'hffffff;
assign target_only_stripe[1426] = 24'hffffff;
assign target_only_stripe[1427] = 24'hffffff;
assign target_only_stripe[1428] = 24'hffffff;
assign target_only_stripe[1429] = 24'hffffff;
assign target_only_stripe[1430] = 24'hffffff;
assign target_only_stripe[1431] = 24'hffffff;
assign target_only_stripe[1432] = 24'hffffff;
assign target_only_stripe[1433] = 24'hffffff;
assign target_only_stripe[1434] = 24'hffffff;
assign target_only_stripe[1435] = 24'hffffff;
assign target_only_stripe[1436] = 24'hffffff;
assign target_only_stripe[1437] = 24'hffffff;
assign target_only_stripe[1438] = 24'hffffff;
assign target_only_stripe[1439] = 24'hffffff;
assign target_only_stripe[1440] = 24'hffffff;
assign target_only_stripe[1441] = 24'hffffff;
assign target_only_stripe[1442] = 24'hffffff;
assign target_only_stripe[1443] = 24'hffffff;
assign target_only_stripe[1444] = 24'hffffff;
assign target_only_stripe[1445] = 24'hffffff;
assign target_only_stripe[1446] = 24'hffffff;
assign target_only_stripe[1447] = 24'hffffff;
assign target_only_stripe[1448] = 24'hffffff;
assign target_only_stripe[1449] = 24'h141414;
assign target_only_stripe[1450] = 24'h000000;
assign target_only_stripe[1451] = 24'h000000;
assign target_only_stripe[1452] = 24'h000000;
assign target_only_stripe[1453] = 24'h000000;
assign target_only_stripe[1454] = 24'h000000;
assign target_only_stripe[1455] = 24'h000000;
assign target_only_stripe[1456] = 24'h000000;
assign target_only_stripe[1457] = 24'h000000;
assign target_only_stripe[1458] = 24'h000000;
assign target_only_stripe[1459] = 24'h000000;
assign target_only_stripe[1460] = 24'h000000;
assign target_only_stripe[1461] = 24'h000000;
assign target_only_stripe[1462] = 24'h000000;
assign target_only_stripe[1463] = 24'h000000;
assign target_only_stripe[1464] = 24'h000000;
assign target_only_stripe[1465] = 24'h000000;
assign target_only_stripe[1466] = 24'h000000;
assign target_only_stripe[1467] = 24'h000000;
assign target_only_stripe[1468] = 24'h000000;
assign target_only_stripe[1469] = 24'h000000;
assign target_only_stripe[1470] = 24'h000000;
assign target_only_stripe[1471] = 24'h000000;
assign target_only_stripe[1472] = 24'h000000;
assign target_only_stripe[1473] = 24'h000000;
assign target_only_stripe[1474] = 24'h000000;
assign target_only_stripe[1475] = 24'h000000;
assign target_only_stripe[1476] = 24'h000000;
assign target_only_stripe[1477] = 24'h000000;
assign target_only_stripe[1478] = 24'h000000;
assign target_only_stripe[1479] = 24'h000000;
assign target_only_stripe[1480] = 24'h000000;
assign target_only_stripe[1481] = 24'h000000;
assign target_only_stripe[1482] = 24'h000000;
assign target_only_stripe[1483] = 24'h000000;
assign target_only_stripe[1484] = 24'h000000;
assign target_only_stripe[1485] = 24'h000000;
assign target_only_stripe[1486] = 24'h000000;
assign target_only_stripe[1487] = 24'h000000;
assign target_only_stripe[1488] = 24'h000000;
assign target_only_stripe[1489] = 24'h000000;
assign target_only_stripe[1490] = 24'h000000;
assign target_only_stripe[1491] = 24'h000000;
assign target_only_stripe[1492] = 24'h000000;
assign target_only_stripe[1493] = 24'h000000;
assign target_only_stripe[1494] = 24'h000000;
assign target_only_stripe[1495] = 24'h000000;
assign target_only_stripe[1496] = 24'h000000;
assign target_only_stripe[1497] = 24'h000000;
assign target_only_stripe[1498] = 24'h000000;
assign target_only_stripe[1499] = 24'h000000;
assign target_only_stripe[1500] = 24'h000000;
assign target_only_stripe[1501] = 24'h000000;
assign target_only_stripe[1502] = 24'h000000;
assign target_only_stripe[1503] = 24'h000000;
assign target_only_stripe[1504] = 24'h000000;
assign target_only_stripe[1505] = 24'h000000;
assign target_only_stripe[1506] = 24'h000000;
assign target_only_stripe[1507] = 24'h000000;
assign target_only_stripe[1508] = 24'h000000;
assign target_only_stripe[1509] = 24'h000000;
assign target_only_stripe[1510] = 24'h000000;
assign target_only_stripe[1511] = 24'h101010;
assign target_only_stripe[1512] = 24'hffffff;
assign target_only_stripe[1513] = 24'hffffff;
assign target_only_stripe[1514] = 24'hffffff;
assign target_only_stripe[1515] = 24'hffffff;
assign target_only_stripe[1516] = 24'hffffff;
assign target_only_stripe[1517] = 24'hffffff;
assign target_only_stripe[1518] = 24'hffffff;
assign target_only_stripe[1519] = 24'hffffff;
assign target_only_stripe[1520] = 24'hffffff;
assign target_only_stripe[1521] = 24'hffffff;
assign target_only_stripe[1522] = 24'hffffff;
assign target_only_stripe[1523] = 24'hffffff;
assign target_only_stripe[1524] = 24'hffffff;
assign target_only_stripe[1525] = 24'hffffff;
assign target_only_stripe[1526] = 24'hffffff;
assign target_only_stripe[1527] = 24'hffffff;
assign target_only_stripe[1528] = 24'hffffff;
assign target_only_stripe[1529] = 24'hffffff;
assign target_only_stripe[1530] = 24'hffffff;
assign target_only_stripe[1531] = 24'hffffff;
assign target_only_stripe[1532] = 24'hffffff;
assign target_only_stripe[1533] = 24'hffffff;
assign target_only_stripe[1534] = 24'hffffff;
assign target_only_stripe[1535] = 24'hffffff;
assign target_only_stripe[1536] = 24'hffffff;
assign target_only_stripe[1537] = 24'hffffff;
assign target_only_stripe[1538] = 24'hffffff;
assign target_only_stripe[1539] = 24'hffffff;
assign target_only_stripe[1540] = 24'hffffff;
assign target_only_stripe[1541] = 24'hffffff;
assign target_only_stripe[1542] = 24'hffffff;
assign target_only_stripe[1543] = 24'hffffff;
assign target_only_stripe[1544] = 24'hffffff;
assign target_only_stripe[1545] = 24'hffffff;
assign target_only_stripe[1546] = 24'h434343;
assign target_only_stripe[1547] = 24'h000000;
assign target_only_stripe[1548] = 24'h000000;
assign target_only_stripe[1549] = 24'h000000;
assign target_only_stripe[1550] = 24'h000000;
assign target_only_stripe[1551] = 24'h000000;
assign target_only_stripe[1552] = 24'h000000;
assign target_only_stripe[1553] = 24'h000000;
assign target_only_stripe[1554] = 24'h000000;
assign target_only_stripe[1555] = 24'h000000;
assign target_only_stripe[1556] = 24'h000000;
assign target_only_stripe[1557] = 24'h000000;
assign target_only_stripe[1558] = 24'h000000;
assign target_only_stripe[1559] = 24'h000000;
assign target_only_stripe[1560] = 24'h000000;
assign target_only_stripe[1561] = 24'h000000;
assign target_only_stripe[1562] = 24'h000000;
assign target_only_stripe[1563] = 24'h000000;
assign target_only_stripe[1564] = 24'h000000;
assign target_only_stripe[1565] = 24'h000000;
assign target_only_stripe[1566] = 24'h000000;
assign target_only_stripe[1567] = 24'h000000;
assign target_only_stripe[1568] = 24'h000000;
assign target_only_stripe[1569] = 24'h000000;
assign target_only_stripe[1570] = 24'h000000;
assign target_only_stripe[1571] = 24'h000000;
assign target_only_stripe[1572] = 24'h000000;
assign target_only_stripe[1573] = 24'h000000;
assign target_only_stripe[1574] = 24'h000000;
assign target_only_stripe[1575] = 24'h000000;
assign target_only_stripe[1576] = 24'h000000;
assign target_only_stripe[1577] = 24'h000000;
assign target_only_stripe[1578] = 24'h0a0a0a;
assign target_only_stripe[1579] = 24'hcecece;
assign target_only_stripe[1580] = 24'hffffff;
assign target_only_stripe[1581] = 24'hfaf7f5;
assign target_only_stripe[1582] = 24'hffffff;
assign target_only_stripe[1583] = 24'hffffff;
assign target_only_stripe[1584] = 24'hffffff;
assign target_only_stripe[1585] = 24'hffffff;
assign target_only_stripe[1586] = 24'hffffff;
assign target_only_stripe[1587] = 24'hffffff;
assign target_only_stripe[1588] = 24'hffffff;
assign target_only_stripe[1589] = 24'hffffff;
assign target_only_stripe[1590] = 24'hffffff;
assign target_only_stripe[1591] = 24'hffffff;
assign target_only_stripe[1592] = 24'hffffff;
assign target_only_stripe[1593] = 24'hffffff;
assign target_only_stripe[1594] = 24'hffffff;
assign target_only_stripe[1595] = 24'hffffff;
assign target_only_stripe[1596] = 24'hffffff;
assign target_only_stripe[1597] = 24'hffffff;
assign target_only_stripe[1598] = 24'hffffff;
assign target_only_stripe[1599] = 24'hffffff;
assign target_only_stripe[1600] = 24'hffffff;
assign target_only_stripe[1601] = 24'hffffff;
assign target_only_stripe[1602] = 24'hffffff;
assign target_only_stripe[1603] = 24'hffffff;
assign target_only_stripe[1604] = 24'hffffff;
assign target_only_stripe[1605] = 24'hffffff;
assign target_only_stripe[1606] = 24'hffffff;
assign target_only_stripe[1607] = 24'hffffff;
assign target_only_stripe[1608] = 24'hffffff;
assign target_only_stripe[1609] = 24'hffffff;
assign target_only_stripe[1610] = 24'hffffff;
assign target_only_stripe[1611] = 24'hffffff;
assign target_only_stripe[1612] = 24'hd2d2d2;
assign target_only_stripe[1613] = 24'h0c0c0c;
assign target_only_stripe[1614] = 24'h000000;
assign target_only_stripe[1615] = 24'h000000;
assign target_only_stripe[1616] = 24'h000000;
assign target_only_stripe[1617] = 24'h000000;
assign target_only_stripe[1618] = 24'h000000;
assign target_only_stripe[1619] = 24'h000000;
assign target_only_stripe[1620] = 24'h000000;
assign target_only_stripe[1621] = 24'h000000;
assign target_only_stripe[1622] = 24'h000000;
assign target_only_stripe[1623] = 24'h000000;
assign target_only_stripe[1624] = 24'h000000;
assign target_only_stripe[1625] = 24'h000000;
assign target_only_stripe[1626] = 24'h000000;
assign target_only_stripe[1627] = 24'h000000;
assign target_only_stripe[1628] = 24'h000000;
assign target_only_stripe[1629] = 24'h000000;
assign target_only_stripe[1630] = 24'h000000;
assign target_only_stripe[1631] = 24'h000000;
assign target_only_stripe[1632] = 24'h000000;
assign target_only_stripe[1633] = 24'h000000;
assign target_only_stripe[1634] = 24'h000000;
assign target_only_stripe[1635] = 24'h000000;
assign target_only_stripe[1636] = 24'h000000;
assign target_only_stripe[1637] = 24'h000000;
assign target_only_stripe[1638] = 24'h000000;
assign target_only_stripe[1639] = 24'h000000;
assign target_only_stripe[1640] = 24'h000000;
assign target_only_stripe[1641] = 24'h000000;
assign target_only_stripe[1642] = 24'h000000;
assign target_only_stripe[1643] = 24'h000000;
assign target_only_stripe[1644] = 24'h000000;
assign target_only_stripe[1645] = 24'h000000;
assign target_only_stripe[1646] = 24'h000000;
assign target_only_stripe[1647] = 24'h000000;
assign target_only_stripe[1648] = 24'h000000;
assign target_only_stripe[1649] = 24'h000000;
assign target_only_stripe[1650] = 24'h000000;
assign target_only_stripe[1651] = 24'h000000;
assign target_only_stripe[1652] = 24'h000000;
assign target_only_stripe[1653] = 24'h000000;
assign target_only_stripe[1654] = 24'h000000;
assign target_only_stripe[1655] = 24'h000000;
assign target_only_stripe[1656] = 24'h000000;
assign target_only_stripe[1657] = 24'h000000;
assign target_only_stripe[1658] = 24'h000000;
assign target_only_stripe[1659] = 24'h000000;
assign target_only_stripe[1660] = 24'h000000;
assign target_only_stripe[1661] = 24'h000000;
assign target_only_stripe[1662] = 24'h000000;
assign target_only_stripe[1663] = 24'h000000;
assign target_only_stripe[1664] = 24'h000000;
assign target_only_stripe[1665] = 24'h000000;
assign target_only_stripe[1666] = 24'h000000;
assign target_only_stripe[1667] = 24'h000000;
assign target_only_stripe[1668] = 24'h000000;
assign target_only_stripe[1669] = 24'h000000;
assign target_only_stripe[1670] = 24'h000000;
assign target_only_stripe[1671] = 24'h000000;
assign target_only_stripe[1672] = 24'h000000;
assign target_only_stripe[1673] = 24'h000000;
assign target_only_stripe[1674] = 24'h000000;
assign target_only_stripe[1675] = 24'h000000;
assign target_only_stripe[1676] = 24'h0c0c0c;
assign target_only_stripe[1677] = 24'hdbdbdb;
assign target_only_stripe[1678] = 24'hffffff;
assign target_only_stripe[1679] = 24'hffffff;
assign target_only_stripe[1680] = 24'hffffff;
assign target_only_stripe[1681] = 24'hffffff;
assign target_only_stripe[1682] = 24'hffffff;
assign target_only_stripe[1683] = 24'hffffff;
assign target_only_stripe[1684] = 24'hffffff;
assign target_only_stripe[1685] = 24'hffffff;
assign target_only_stripe[1686] = 24'hffffff;
assign target_only_stripe[1687] = 24'hffffff;
assign target_only_stripe[1688] = 24'hffffff;
assign target_only_stripe[1689] = 24'hffffff;
assign target_only_stripe[1690] = 24'hffffff;
assign target_only_stripe[1691] = 24'hffffff;
assign target_only_stripe[1692] = 24'hffffff;
assign target_only_stripe[1693] = 24'hffffff;
assign target_only_stripe[1694] = 24'hffffff;
assign target_only_stripe[1695] = 24'hffffff;
assign target_only_stripe[1696] = 24'hffffff;
assign target_only_stripe[1697] = 24'hffffff;
assign target_only_stripe[1698] = 24'hffffff;
assign target_only_stripe[1699] = 24'hffffff;
assign target_only_stripe[1700] = 24'hffffff;
assign target_only_stripe[1701] = 24'hffffff;
assign target_only_stripe[1702] = 24'hffffff;
assign target_only_stripe[1703] = 24'hffffff;
assign target_only_stripe[1704] = 24'hffffff;
assign target_only_stripe[1705] = 24'hffffff;
assign target_only_stripe[1706] = 24'hffffff;
assign target_only_stripe[1707] = 24'hffffff;
assign target_only_stripe[1708] = 24'hffffff;
assign target_only_stripe[1709] = 24'hffffff;
assign target_only_stripe[1710] = 24'hcdcdcd;
assign target_only_stripe[1711] = 24'h050505;
assign target_only_stripe[1712] = 24'h000000;
assign target_only_stripe[1713] = 24'h000000;
assign target_only_stripe[1714] = 24'h000000;
assign target_only_stripe[1715] = 24'h000000;
assign target_only_stripe[1716] = 24'h000000;
assign target_only_stripe[1717] = 24'h000000;
assign target_only_stripe[1718] = 24'h000000;
assign target_only_stripe[1719] = 24'h000000;
assign target_only_stripe[1720] = 24'h000000;
assign target_only_stripe[1721] = 24'h000000;
assign target_only_stripe[1722] = 24'h000000;
assign target_only_stripe[1723] = 24'h000000;
assign target_only_stripe[1724] = 24'h000000;
assign target_only_stripe[1725] = 24'h000000;
assign target_only_stripe[1726] = 24'h000000;
assign target_only_stripe[1727] = 24'h000000;
assign target_only_stripe[1728] = 24'h000000;
assign target_only_stripe[1729] = 24'h000000;
assign target_only_stripe[1730] = 24'h000000;
assign target_only_stripe[1731] = 24'h000000;
assign target_only_stripe[1732] = 24'h000000;
assign target_only_stripe[1733] = 24'h000000;
assign target_only_stripe[1734] = 24'h000000;
assign target_only_stripe[1735] = 24'h000000;
assign target_only_stripe[1736] = 24'h000000;
assign target_only_stripe[1737] = 24'h000000;
assign target_only_stripe[1738] = 24'h000000;
assign target_only_stripe[1739] = 24'h000000;
assign target_only_stripe[1740] = 24'h000000;
assign target_only_stripe[1741] = 24'h000000;
assign target_only_stripe[1742] = 24'h000000;
assign target_only_stripe[1743] = 24'hf2f2f2;
assign target_only_stripe[1744] = 24'hffffff;
assign target_only_stripe[1745] = 24'hffffff;
assign target_only_stripe[1746] = 24'hffffff;
assign target_only_stripe[1747] = 24'hffffff;
assign target_only_stripe[1748] = 24'hffffff;
assign target_only_stripe[1749] = 24'hffffff;
assign target_only_stripe[1750] = 24'hffffff;
assign target_only_stripe[1751] = 24'hffffff;
assign target_only_stripe[1752] = 24'hffffff;
assign target_only_stripe[1753] = 24'hffffff;
assign target_only_stripe[1754] = 24'hffffff;
assign target_only_stripe[1755] = 24'hffffff;
assign target_only_stripe[1756] = 24'hffffff;
assign target_only_stripe[1757] = 24'hffffff;
assign target_only_stripe[1758] = 24'hffffff;
assign target_only_stripe[1759] = 24'hffffff;
assign target_only_stripe[1760] = 24'hffffff;
assign target_only_stripe[1761] = 24'hffffff;
assign target_only_stripe[1762] = 24'hffffff;
assign target_only_stripe[1763] = 24'hffffff;
assign target_only_stripe[1764] = 24'hffffff;
assign target_only_stripe[1765] = 24'hffffff;
assign target_only_stripe[1766] = 24'hffffff;
assign target_only_stripe[1767] = 24'hffffff;
assign target_only_stripe[1768] = 24'hffffff;
assign target_only_stripe[1769] = 24'hffffff;
assign target_only_stripe[1770] = 24'hffffff;
assign target_only_stripe[1771] = 24'hffffff;
assign target_only_stripe[1772] = 24'hffffff;
assign target_only_stripe[1773] = 24'hffffff;
assign target_only_stripe[1774] = 24'hffffff;
assign target_only_stripe[1775] = 24'hffffff;
assign target_only_stripe[1776] = 24'hffffff;
assign target_only_stripe[1777] = 24'hb4b4b4;
assign target_only_stripe[1778] = 24'h000000;
assign target_only_stripe[1779] = 24'h000000;
assign target_only_stripe[1780] = 24'h000000;
assign target_only_stripe[1781] = 24'h000000;
assign target_only_stripe[1782] = 24'h000000;
assign target_only_stripe[1783] = 24'h000000;
assign target_only_stripe[1784] = 24'h000000;
assign target_only_stripe[1785] = 24'h000000;
assign target_only_stripe[1786] = 24'h000000;
assign target_only_stripe[1787] = 24'h000000;
assign target_only_stripe[1788] = 24'h000000;
assign target_only_stripe[1789] = 24'h000000;
assign target_only_stripe[1790] = 24'h000000;
assign target_only_stripe[1791] = 24'h000000;
assign target_only_stripe[1792] = 24'h000000;
assign target_only_stripe[1793] = 24'h000000;
assign target_only_stripe[1794] = 24'h000000;
assign target_only_stripe[1795] = 24'h000000;
assign target_only_stripe[1796] = 24'h000000;
assign target_only_stripe[1797] = 24'h000000;
assign target_only_stripe[1798] = 24'h000000;
assign target_only_stripe[1799] = 24'h000000;
assign target_only_stripe[1800] = 24'h000000;
assign target_only_stripe[1801] = 24'h000000;
assign target_only_stripe[1802] = 24'h000000;
assign target_only_stripe[1803] = 24'h000000;
assign target_only_stripe[1804] = 24'h000000;
assign target_only_stripe[1805] = 24'h000000;
assign target_only_stripe[1806] = 24'h000000;
assign target_only_stripe[1807] = 24'h000000;
assign target_only_stripe[1808] = 24'h000000;
assign target_only_stripe[1809] = 24'h000000;
assign target_only_stripe[1810] = 24'h000000;
assign target_only_stripe[1811] = 24'h000000;
assign target_only_stripe[1812] = 24'h000000;
assign target_only_stripe[1813] = 24'h000000;
assign target_only_stripe[1814] = 24'h000000;
assign target_only_stripe[1815] = 24'h000000;
assign target_only_stripe[1816] = 24'h000000;
assign target_only_stripe[1817] = 24'h000000;
assign target_only_stripe[1818] = 24'h000000;
assign target_only_stripe[1819] = 24'h000000;
assign target_only_stripe[1820] = 24'h000000;
assign target_only_stripe[1821] = 24'h000000;
assign target_only_stripe[1822] = 24'h000000;
assign target_only_stripe[1823] = 24'h000000;
assign target_only_stripe[1824] = 24'h000000;
assign target_only_stripe[1825] = 24'h000000;
assign target_only_stripe[1826] = 24'h000000;
assign target_only_stripe[1827] = 24'h000000;
assign target_only_stripe[1828] = 24'h000000;
assign target_only_stripe[1829] = 24'h000000;
assign target_only_stripe[1830] = 24'h000000;
assign target_only_stripe[1831] = 24'h000000;
assign target_only_stripe[1832] = 24'h000000;
assign target_only_stripe[1833] = 24'h000000;
assign target_only_stripe[1834] = 24'h000000;
assign target_only_stripe[1835] = 24'h000000;
assign target_only_stripe[1836] = 24'h000000;
assign target_only_stripe[1837] = 24'h000000;
assign target_only_stripe[1838] = 24'h000000;
assign target_only_stripe[1839] = 24'h000000;
assign target_only_stripe[1840] = 24'h000000;
assign target_only_stripe[1841] = 24'hacacac;
assign target_only_stripe[1842] = 24'hffffff;
assign target_only_stripe[1843] = 24'hffffff;
assign target_only_stripe[1844] = 24'hffffff;
assign target_only_stripe[1845] = 24'hffffff;
assign target_only_stripe[1846] = 24'hffffff;
assign target_only_stripe[1847] = 24'hffffff;
assign target_only_stripe[1848] = 24'hffffff;
assign target_only_stripe[1849] = 24'hffffff;
assign target_only_stripe[1850] = 24'hffffff;
assign target_only_stripe[1851] = 24'hffffff;
assign target_only_stripe[1852] = 24'hffffff;
assign target_only_stripe[1853] = 24'hffffff;
assign target_only_stripe[1854] = 24'hffffff;
assign target_only_stripe[1855] = 24'hffffff;
assign target_only_stripe[1856] = 24'hffffff;
assign target_only_stripe[1857] = 24'hffffff;
assign target_only_stripe[1858] = 24'hffffff;
assign target_only_stripe[1859] = 24'hffffff;
assign target_only_stripe[1860] = 24'hffffff;
assign target_only_stripe[1861] = 24'hffffff;
assign target_only_stripe[1862] = 24'hffffff;
assign target_only_stripe[1863] = 24'hffffff;
assign target_only_stripe[1864] = 24'hffffff;
assign target_only_stripe[1865] = 24'hffffff;
assign target_only_stripe[1866] = 24'hffffff;
assign target_only_stripe[1867] = 24'hffffff;
assign target_only_stripe[1868] = 24'hffffff;
assign target_only_stripe[1869] = 24'hffffff;
assign target_only_stripe[1870] = 24'hffffff;
assign target_only_stripe[1871] = 24'hffffff;
assign target_only_stripe[1872] = 24'hffffff;
assign target_only_stripe[1873] = 24'hffffff;
assign target_only_stripe[1874] = 24'hffffff;
assign target_only_stripe[1875] = 24'hffffff;
assign target_only_stripe[1876] = 24'h000000;
assign target_only_stripe[1877] = 24'h000000;
assign target_only_stripe[1878] = 24'h000000;
assign target_only_stripe[1879] = 24'h000000;
assign target_only_stripe[1880] = 24'h000000;
assign target_only_stripe[1881] = 24'h000000;
assign target_only_stripe[1882] = 24'h000000;
assign target_only_stripe[1883] = 24'h000000;
assign target_only_stripe[1884] = 24'h000000;
assign target_only_stripe[1885] = 24'h000000;
assign target_only_stripe[1886] = 24'h000000;
assign target_only_stripe[1887] = 24'h000000;
assign target_only_stripe[1888] = 24'h000000;
assign target_only_stripe[1889] = 24'h000000;
assign target_only_stripe[1890] = 24'h000000;
assign target_only_stripe[1891] = 24'h000000;
assign target_only_stripe[1892] = 24'h000000;
assign target_only_stripe[1893] = 24'h000000;
assign target_only_stripe[1894] = 24'h000000;
assign target_only_stripe[1895] = 24'h000000;
assign target_only_stripe[1896] = 24'h000000;
assign target_only_stripe[1897] = 24'h000000;
assign target_only_stripe[1898] = 24'h000000;
assign target_only_stripe[1899] = 24'h000000;
assign target_only_stripe[1900] = 24'h000000;
assign target_only_stripe[1901] = 24'h000000;
assign target_only_stripe[1902] = 24'h000000;
assign target_only_stripe[1903] = 24'h000000;
assign target_only_stripe[1904] = 24'h000000;
assign target_only_stripe[1905] = 24'h000000;
assign target_only_stripe[1906] = 24'h000000;
assign target_only_stripe[1907] = 24'h030303;
assign target_only_stripe[1908] = 24'hc7c7c7;
assign target_only_stripe[1909] = 24'hffffff;
assign target_only_stripe[1910] = 24'hffffff;
assign target_only_stripe[1911] = 24'hffffff;
assign target_only_stripe[1912] = 24'hffffff;
assign target_only_stripe[1913] = 24'hffffff;
assign target_only_stripe[1914] = 24'hffffff;
assign target_only_stripe[1915] = 24'hffffff;
assign target_only_stripe[1916] = 24'hffffff;
assign target_only_stripe[1917] = 24'hffffff;
assign target_only_stripe[1918] = 24'hffffff;
assign target_only_stripe[1919] = 24'hffffff;
assign target_only_stripe[1920] = 24'hffffff;
assign target_only_stripe[1921] = 24'hffffff;
assign target_only_stripe[1922] = 24'hffffff;
assign target_only_stripe[1923] = 24'hffffff;
assign target_only_stripe[1924] = 24'hffffff;
assign target_only_stripe[1925] = 24'hffffff;
assign target_only_stripe[1926] = 24'hffffff;
assign target_only_stripe[1927] = 24'hffffff;
assign target_only_stripe[1928] = 24'hffffff;
assign target_only_stripe[1929] = 24'hffffff;
assign target_only_stripe[1930] = 24'hffffff;
assign target_only_stripe[1931] = 24'hffffff;
assign target_only_stripe[1932] = 24'hffffff;
assign target_only_stripe[1933] = 24'hffffff;
assign target_only_stripe[1934] = 24'hffffff;
assign target_only_stripe[1935] = 24'hffffff;
assign target_only_stripe[1936] = 24'hffffff;
assign target_only_stripe[1937] = 24'hffffff;
assign target_only_stripe[1938] = 24'hffffff;
assign target_only_stripe[1939] = 24'hffffff;
assign target_only_stripe[1940] = 24'hffffff;
assign target_only_stripe[1941] = 24'hdfdfdf;
assign target_only_stripe[1942] = 24'h141414;
assign target_only_stripe[1943] = 24'h000000;
assign target_only_stripe[1944] = 24'h000000;
assign target_only_stripe[1945] = 24'h000000;
assign target_only_stripe[1946] = 24'h000000;
assign target_only_stripe[1947] = 24'h000000;
assign target_only_stripe[1948] = 24'h000000;
assign target_only_stripe[1949] = 24'h000000;
assign target_only_stripe[1950] = 24'h000000;
assign target_only_stripe[1951] = 24'h000000;
assign target_only_stripe[1952] = 24'h000000;
assign target_only_stripe[1953] = 24'h000000;
assign target_only_stripe[1954] = 24'h000000;
assign target_only_stripe[1955] = 24'h000000;
assign target_only_stripe[1956] = 24'h000000;
assign target_only_stripe[1957] = 24'h000000;
assign target_only_stripe[1958] = 24'h000000;
assign target_only_stripe[1959] = 24'h000000;
assign target_only_stripe[1960] = 24'h000000;
assign target_only_stripe[1961] = 24'h000000;
assign target_only_stripe[1962] = 24'h000000;
assign target_only_stripe[1963] = 24'h000000;
assign target_only_stripe[1964] = 24'h000000;
assign target_only_stripe[1965] = 24'h000000;
assign target_only_stripe[1966] = 24'h000000;
assign target_only_stripe[1967] = 24'h000000;
assign target_only_stripe[1968] = 24'h000000;
assign target_only_stripe[1969] = 24'h000000;
assign target_only_stripe[1970] = 24'h000000;
assign target_only_stripe[1971] = 24'h000000;
assign target_only_stripe[1972] = 24'h000000;
assign target_only_stripe[1973] = 24'h000000;
assign target_only_stripe[1974] = 24'h000000;
assign target_only_stripe[1975] = 24'h000000;
assign target_only_stripe[1976] = 24'h000000;
assign target_only_stripe[1977] = 24'h000000;
assign target_only_stripe[1978] = 24'h000000;
assign target_only_stripe[1979] = 24'h000000;
assign target_only_stripe[1980] = 24'h000000;
assign target_only_stripe[1981] = 24'h000000;
assign target_only_stripe[1982] = 24'h000000;
assign target_only_stripe[1983] = 24'h000000;
assign target_only_stripe[1984] = 24'h000000;
assign target_only_stripe[1985] = 24'h000000;
assign target_only_stripe[1986] = 24'h000000;
assign target_only_stripe[1987] = 24'h000000;
assign target_only_stripe[1988] = 24'h000000;
assign target_only_stripe[1989] = 24'h000000;
assign target_only_stripe[1990] = 24'h000000;
assign target_only_stripe[1991] = 24'h000000;
assign target_only_stripe[1992] = 24'h000000;
assign target_only_stripe[1993] = 24'h000000;
assign target_only_stripe[1994] = 24'h000000;
assign target_only_stripe[1995] = 24'h000000;
assign target_only_stripe[1996] = 24'h000000;
assign target_only_stripe[1997] = 24'h000000;
assign target_only_stripe[1998] = 24'h000000;
assign target_only_stripe[1999] = 24'h000000;
assign target_only_stripe[2000] = 24'h000000;
assign target_only_stripe[2001] = 24'h000000;
assign target_only_stripe[2002] = 24'h000000;
assign target_only_stripe[2003] = 24'h000000;
assign target_only_stripe[2004] = 24'h000000;
assign target_only_stripe[2005] = 24'h101010;
assign target_only_stripe[2006] = 24'he4e4e4;
assign target_only_stripe[2007] = 24'hffffff;
assign target_only_stripe[2008] = 24'hffffff;
assign target_only_stripe[2009] = 24'hffffff;
assign target_only_stripe[2010] = 24'hffffff;
assign target_only_stripe[2011] = 24'hffffff;
assign target_only_stripe[2012] = 24'hffffff;
assign target_only_stripe[2013] = 24'hffffff;
assign target_only_stripe[2014] = 24'hffffff;
assign target_only_stripe[2015] = 24'hffffff;
assign target_only_stripe[2016] = 24'hffffff;
assign target_only_stripe[2017] = 24'hffffff;
assign target_only_stripe[2018] = 24'hffffff;
assign target_only_stripe[2019] = 24'hffffff;
assign target_only_stripe[2020] = 24'hffffff;
assign target_only_stripe[2021] = 24'hffffff;
assign target_only_stripe[2022] = 24'hffffff;
assign target_only_stripe[2023] = 24'hffffff;
assign target_only_stripe[2024] = 24'hffffff;
assign target_only_stripe[2025] = 24'hffffff;
assign target_only_stripe[2026] = 24'hffffff;
assign target_only_stripe[2027] = 24'hffffff;
assign target_only_stripe[2028] = 24'hffffff;
assign target_only_stripe[2029] = 24'hffffff;
assign target_only_stripe[2030] = 24'hffffff;
assign target_only_stripe[2031] = 24'hffffff;
assign target_only_stripe[2032] = 24'hffffff;
assign target_only_stripe[2033] = 24'hffffff;
assign target_only_stripe[2034] = 24'hffffff;
assign target_only_stripe[2035] = 24'hffffff;
assign target_only_stripe[2036] = 24'hffffff;
assign target_only_stripe[2037] = 24'hffffff;
assign target_only_stripe[2038] = 24'hffffff;
assign target_only_stripe[2039] = 24'hcacaca;
assign target_only_stripe[2040] = 24'h000000;
assign target_only_stripe[2041] = 24'h000000;
assign target_only_stripe[2042] = 24'h000000;
assign target_only_stripe[2043] = 24'h000000;
assign target_only_stripe[2044] = 24'h000000;
assign target_only_stripe[2045] = 24'h000000;
assign target_only_stripe[2046] = 24'h000000;
assign target_only_stripe[2047] = 24'h000000;
assign target_only_stripe[2048] = 24'h000000;
assign target_only_stripe[2049] = 24'h000000;
assign target_only_stripe[2050] = 24'h000000;
assign target_only_stripe[2051] = 24'h000000;
assign target_only_stripe[2052] = 24'h000000;
assign target_only_stripe[2053] = 24'h000000;
assign target_only_stripe[2054] = 24'h000000;
assign target_only_stripe[2055] = 24'h000000;
assign target_only_stripe[2056] = 24'h000000;
assign target_only_stripe[2057] = 24'h000000;
assign target_only_stripe[2058] = 24'h000000;
assign target_only_stripe[2059] = 24'h000000;
assign target_only_stripe[2060] = 24'h000000;
assign target_only_stripe[2061] = 24'h000000;
assign target_only_stripe[2062] = 24'h000000;
assign target_only_stripe[2063] = 24'h000000;
assign target_only_stripe[2064] = 24'h000000;
assign target_only_stripe[2065] = 24'h000000;
assign target_only_stripe[2066] = 24'h000000;
assign target_only_stripe[2067] = 24'h000000;
assign target_only_stripe[2068] = 24'h000000;
assign target_only_stripe[2069] = 24'h000000;
assign target_only_stripe[2070] = 24'h000000;
assign target_only_stripe[2071] = 24'h000000;
assign target_only_stripe[2072] = 24'hffffff;
assign target_only_stripe[2073] = 24'hffffff;
assign target_only_stripe[2074] = 24'hffffff;
assign target_only_stripe[2075] = 24'hffffff;
assign target_only_stripe[2076] = 24'hffffff;
assign target_only_stripe[2077] = 24'hffffff;
assign target_only_stripe[2078] = 24'hffffff;
assign target_only_stripe[2079] = 24'hffffff;
assign target_only_stripe[2080] = 24'hffffff;
assign target_only_stripe[2081] = 24'hffffff;
assign target_only_stripe[2082] = 24'hffffff;
assign target_only_stripe[2083] = 24'hffffff;
assign target_only_stripe[2084] = 24'hffffff;
assign target_only_stripe[2085] = 24'hffffff;
assign target_only_stripe[2086] = 24'hffffff;
assign target_only_stripe[2087] = 24'hffffff;
assign target_only_stripe[2088] = 24'hffffff;
assign target_only_stripe[2089] = 24'hffffff;
assign target_only_stripe[2090] = 24'hffffff;
assign target_only_stripe[2091] = 24'hffffff;
assign target_only_stripe[2092] = 24'hffffff;
assign target_only_stripe[2093] = 24'hffffff;
assign target_only_stripe[2094] = 24'hffffff;
assign target_only_stripe[2095] = 24'hffffff;
assign target_only_stripe[2096] = 24'hffffff;
assign target_only_stripe[2097] = 24'hffffff;
assign target_only_stripe[2098] = 24'hffffff;
assign target_only_stripe[2099] = 24'hffffff;
assign target_only_stripe[2100] = 24'hffffff;
assign target_only_stripe[2101] = 24'hffffff;
assign target_only_stripe[2102] = 24'hffffff;
assign target_only_stripe[2103] = 24'hffffff;
assign target_only_stripe[2104] = 24'hffffff;
assign target_only_stripe[2105] = 24'hffffff;
assign target_only_stripe[2106] = 24'h929292;
assign target_only_stripe[2107] = 24'h000000;
assign target_only_stripe[2108] = 24'h000000;
assign target_only_stripe[2109] = 24'h000000;
assign target_only_stripe[2110] = 24'h000000;
assign target_only_stripe[2111] = 24'h000000;
assign target_only_stripe[2112] = 24'h000000;
assign target_only_stripe[2113] = 24'h000000;
assign target_only_stripe[2114] = 24'h000000;
assign target_only_stripe[2115] = 24'h000000;
assign target_only_stripe[2116] = 24'h000000;
assign target_only_stripe[2117] = 24'h000000;
assign target_only_stripe[2118] = 24'h000000;
assign target_only_stripe[2119] = 24'h000000;
assign target_only_stripe[2120] = 24'h000000;
assign target_only_stripe[2121] = 24'h000000;
assign target_only_stripe[2122] = 24'h000000;
assign target_only_stripe[2123] = 24'h000000;
assign target_only_stripe[2124] = 24'h000000;
assign target_only_stripe[2125] = 24'h000000;
assign target_only_stripe[2126] = 24'h000000;
assign target_only_stripe[2127] = 24'h000000;
assign target_only_stripe[2128] = 24'h000000;
assign target_only_stripe[2129] = 24'h000000;
assign target_only_stripe[2130] = 24'h000000;
assign target_only_stripe[2131] = 24'h000000;
assign target_only_stripe[2132] = 24'h000000;
assign target_only_stripe[2133] = 24'h000000;
assign target_only_stripe[2134] = 24'h000000;
assign target_only_stripe[2135] = 24'h000000;
assign target_only_stripe[2136] = 24'h000000;
assign target_only_stripe[2137] = 24'h000000;
assign target_only_stripe[2138] = 24'h000000;
assign target_only_stripe[2139] = 24'h000000;
assign target_only_stripe[2140] = 24'h000000;
assign target_only_stripe[2141] = 24'h000000;
assign target_only_stripe[2142] = 24'h000000;
assign target_only_stripe[2143] = 24'h000000;
assign target_only_stripe[2144] = 24'h000000;
assign target_only_stripe[2145] = 24'h000000;
assign target_only_stripe[2146] = 24'h000000;
assign target_only_stripe[2147] = 24'h000000;
assign target_only_stripe[2148] = 24'h000000;
assign target_only_stripe[2149] = 24'h000000;
assign target_only_stripe[2150] = 24'h000000;
assign target_only_stripe[2151] = 24'h000000;
assign target_only_stripe[2152] = 24'h000000;
assign target_only_stripe[2153] = 24'h000000;
assign target_only_stripe[2154] = 24'h000000;
assign target_only_stripe[2155] = 24'h000000;
assign target_only_stripe[2156] = 24'h000000;
assign target_only_stripe[2157] = 24'h000000;
assign target_only_stripe[2158] = 24'h000000;
assign target_only_stripe[2159] = 24'h000000;
assign target_only_stripe[2160] = 24'h000000;
assign target_only_stripe[2161] = 24'h000000;
assign target_only_stripe[2162] = 24'h000000;
assign target_only_stripe[2163] = 24'h000000;
assign target_only_stripe[2164] = 24'h000000;
assign target_only_stripe[2165] = 24'h000000;
assign target_only_stripe[2166] = 24'h000000;
assign target_only_stripe[2167] = 24'h000000;
assign target_only_stripe[2168] = 24'h000000;
assign target_only_stripe[2169] = 24'h000000;
assign target_only_stripe[2170] = 24'h959595;
assign target_only_stripe[2171] = 24'hffffff;
assign target_only_stripe[2172] = 24'hffffff;
assign target_only_stripe[2173] = 24'hffffff;
assign target_only_stripe[2174] = 24'hffffff;
assign target_only_stripe[2175] = 24'hffffff;
assign target_only_stripe[2176] = 24'hffffff;
assign target_only_stripe[2177] = 24'hffffff;
assign target_only_stripe[2178] = 24'hffffff;
assign target_only_stripe[2179] = 24'hffffff;
assign target_only_stripe[2180] = 24'hffffff;
assign target_only_stripe[2181] = 24'hffffff;
assign target_only_stripe[2182] = 24'hffffff;
assign target_only_stripe[2183] = 24'hffffff;
assign target_only_stripe[2184] = 24'hffffff;
assign target_only_stripe[2185] = 24'hffffff;
assign target_only_stripe[2186] = 24'hffffff;
assign target_only_stripe[2187] = 24'hffffff;
assign target_only_stripe[2188] = 24'hffffff;
assign target_only_stripe[2189] = 24'hffffff;
assign target_only_stripe[2190] = 24'hffffff;
assign target_only_stripe[2191] = 24'hffffff;
assign target_only_stripe[2192] = 24'hffffff;
assign target_only_stripe[2193] = 24'hffffff;
assign target_only_stripe[2194] = 24'hffffff;
assign target_only_stripe[2195] = 24'hffffff;
assign target_only_stripe[2196] = 24'hffffff;
assign target_only_stripe[2197] = 24'hffffff;
assign target_only_stripe[2198] = 24'hffffff;
assign target_only_stripe[2199] = 24'hffffff;
assign target_only_stripe[2200] = 24'hffffff;
assign target_only_stripe[2201] = 24'hffffff;
assign target_only_stripe[2202] = 24'hffffff;
assign target_only_stripe[2203] = 24'hffffff;
assign target_only_stripe[2204] = 24'hffffff;
assign target_only_stripe[2205] = 24'h000000;
assign target_only_stripe[2206] = 24'h000000;
assign target_only_stripe[2207] = 24'h000000;
assign target_only_stripe[2208] = 24'h000000;
assign target_only_stripe[2209] = 24'h000000;
assign target_only_stripe[2210] = 24'h000000;
assign target_only_stripe[2211] = 24'h000000;
assign target_only_stripe[2212] = 24'h000000;
assign target_only_stripe[2213] = 24'h000000;
assign target_only_stripe[2214] = 24'h000000;
assign target_only_stripe[2215] = 24'h000000;
assign target_only_stripe[2216] = 24'h000000;
assign target_only_stripe[2217] = 24'h000000;
assign target_only_stripe[2218] = 24'h000000;
assign target_only_stripe[2219] = 24'h000000;
assign target_only_stripe[2220] = 24'h000000;
assign target_only_stripe[2221] = 24'h000000;
assign target_only_stripe[2222] = 24'h000000;
assign target_only_stripe[2223] = 24'h000000;
assign target_only_stripe[2224] = 24'h000000;
assign target_only_stripe[2225] = 24'h000000;
assign target_only_stripe[2226] = 24'h000000;
assign target_only_stripe[2227] = 24'h000000;
assign target_only_stripe[2228] = 24'h000000;
assign target_only_stripe[2229] = 24'h000000;
assign target_only_stripe[2230] = 24'h000000;
assign target_only_stripe[2231] = 24'h000000;
assign target_only_stripe[2232] = 24'h000000;
assign target_only_stripe[2233] = 24'h000000;
assign target_only_stripe[2234] = 24'h000000;
assign target_only_stripe[2235] = 24'h000000;
assign target_only_stripe[2236] = 24'h000000;
assign target_only_stripe[2237] = 24'hc4c4c4;
assign target_only_stripe[2238] = 24'hffffff;
assign target_only_stripe[2239] = 24'hffffff;
assign target_only_stripe[2240] = 24'hffffff;
assign target_only_stripe[2241] = 24'hffffff;
assign target_only_stripe[2242] = 24'hffffff;
assign target_only_stripe[2243] = 24'hffffff;
assign target_only_stripe[2244] = 24'hffffff;
assign target_only_stripe[2245] = 24'hffffff;
assign target_only_stripe[2246] = 24'hffffff;
assign target_only_stripe[2247] = 24'hffffff;
assign target_only_stripe[2248] = 24'hffffff;
assign target_only_stripe[2249] = 24'hffffff;
assign target_only_stripe[2250] = 24'hffffff;
assign target_only_stripe[2251] = 24'hffffff;
assign target_only_stripe[2252] = 24'hffffff;
assign target_only_stripe[2253] = 24'hffffff;
assign target_only_stripe[2254] = 24'hffffff;
assign target_only_stripe[2255] = 24'hffffff;
assign target_only_stripe[2256] = 24'hffffff;
assign target_only_stripe[2257] = 24'hffffff;
assign target_only_stripe[2258] = 24'hffffff;
assign target_only_stripe[2259] = 24'hffffff;
assign target_only_stripe[2260] = 24'hffffff;
assign target_only_stripe[2261] = 24'hffffff;
assign target_only_stripe[2262] = 24'hffffff;
assign target_only_stripe[2263] = 24'hffffff;
assign target_only_stripe[2264] = 24'hffffff;
assign target_only_stripe[2265] = 24'hffffff;
assign target_only_stripe[2266] = 24'hffffff;
assign target_only_stripe[2267] = 24'hffffff;
assign target_only_stripe[2268] = 24'hffffff;
assign target_only_stripe[2269] = 24'hffffff;
assign target_only_stripe[2270] = 24'he8e8e8;
assign target_only_stripe[2271] = 24'h181818;
assign target_only_stripe[2272] = 24'h000000;
assign target_only_stripe[2273] = 24'h000000;
assign target_only_stripe[2274] = 24'h000000;
assign target_only_stripe[2275] = 24'h000000;
assign target_only_stripe[2276] = 24'h000000;
assign target_only_stripe[2277] = 24'h000000;
assign target_only_stripe[2278] = 24'h000000;
assign target_only_stripe[2279] = 24'h000000;
assign target_only_stripe[2280] = 24'h000000;
assign target_only_stripe[2281] = 24'h000000;
assign target_only_stripe[2282] = 24'h000000;
assign target_only_stripe[2283] = 24'h000000;
assign target_only_stripe[2284] = 24'h000000;
assign target_only_stripe[2285] = 24'h000000;
assign target_only_stripe[2286] = 24'h000000;
assign target_only_stripe[2287] = 24'h000000;
assign target_only_stripe[2288] = 24'h000000;
assign target_only_stripe[2289] = 24'h000000;
assign target_only_stripe[2290] = 24'h000000;
assign target_only_stripe[2291] = 24'h000000;
assign target_only_stripe[2292] = 24'h000000;
assign target_only_stripe[2293] = 24'h000000;
assign target_only_stripe[2294] = 24'h000000;
assign target_only_stripe[2295] = 24'h000000;
assign target_only_stripe[2296] = 24'h000000;
assign target_only_stripe[2297] = 24'h000000;
assign target_only_stripe[2298] = 24'h000000;
assign target_only_stripe[2299] = 24'h000000;
assign target_only_stripe[2300] = 24'h000000;
assign target_only_stripe[2301] = 24'h000000;
assign target_only_stripe[2302] = 24'h000000;
assign target_only_stripe[2303] = 24'h000000;
assign target_only_stripe[2304] = 24'h000000;
assign target_only_stripe[2305] = 24'h000000;
assign target_only_stripe[2306] = 24'h000000;
assign target_only_stripe[2307] = 24'h000000;
assign target_only_stripe[2308] = 24'h000000;
assign target_only_stripe[2309] = 24'h000000;
assign target_only_stripe[2310] = 24'h000000;
assign target_only_stripe[2311] = 24'h000000;
assign target_only_stripe[2312] = 24'h000000;
assign target_only_stripe[2313] = 24'h000000;
assign target_only_stripe[2314] = 24'h000000;
assign target_only_stripe[2315] = 24'h000000;
assign target_only_stripe[2316] = 24'h000000;
assign target_only_stripe[2317] = 24'h000000;
assign target_only_stripe[2318] = 24'h000000;
assign target_only_stripe[2319] = 24'h000000;
assign target_only_stripe[2320] = 24'h000000;
assign target_only_stripe[2321] = 24'h000000;
assign target_only_stripe[2322] = 24'h000000;
assign target_only_stripe[2323] = 24'h000000;
assign target_only_stripe[2324] = 24'h000000;
assign target_only_stripe[2325] = 24'h000000;
assign target_only_stripe[2326] = 24'h000000;
assign target_only_stripe[2327] = 24'h000000;
assign target_only_stripe[2328] = 24'h000000;
assign target_only_stripe[2329] = 24'h000000;
assign target_only_stripe[2330] = 24'h000000;
assign target_only_stripe[2331] = 24'h000000;
assign target_only_stripe[2332] = 24'h000000;
assign target_only_stripe[2333] = 24'h000000;
assign target_only_stripe[2334] = 24'h111111;
assign target_only_stripe[2335] = 24'he8e8e8;
assign target_only_stripe[2336] = 24'hffffff;
assign target_only_stripe[2337] = 24'hffffff;
assign target_only_stripe[2338] = 24'hffffff;
assign target_only_stripe[2339] = 24'hffffff;
assign target_only_stripe[2340] = 24'hffffff;
assign target_only_stripe[2341] = 24'hffffff;
assign target_only_stripe[2342] = 24'hffffff;
assign target_only_stripe[2343] = 24'hffffff;
assign target_only_stripe[2344] = 24'hffffff;
assign target_only_stripe[2345] = 24'hffffff;
assign target_only_stripe[2346] = 24'hffffff;
assign target_only_stripe[2347] = 24'hffffff;
assign target_only_stripe[2348] = 24'hffffff;
assign target_only_stripe[2349] = 24'hffffff;
assign target_only_stripe[2350] = 24'hffffff;
assign target_only_stripe[2351] = 24'hffffff;
assign target_only_stripe[2352] = 24'hffffff;
assign target_only_stripe[2353] = 24'hffffff;
assign target_only_stripe[2354] = 24'hffffff;
assign target_only_stripe[2355] = 24'hffffff;
assign target_only_stripe[2356] = 24'hffffff;
assign target_only_stripe[2357] = 24'hffffff;
assign target_only_stripe[2358] = 24'hffffff;
assign target_only_stripe[2359] = 24'hffffff;
assign target_only_stripe[2360] = 24'hffffff;
assign target_only_stripe[2361] = 24'hffffff;
assign target_only_stripe[2362] = 24'hffffff;
assign target_only_stripe[2363] = 24'hffffff;
assign target_only_stripe[2364] = 24'hffffff;
assign target_only_stripe[2365] = 24'hffffff;
assign target_only_stripe[2366] = 24'hffffff;
assign target_only_stripe[2367] = 24'hffffff;
assign target_only_stripe[2368] = 24'hbebebe;
assign target_only_stripe[2369] = 24'h000000;
assign target_only_stripe[2370] = 24'h000000;
assign target_only_stripe[2371] = 24'h000000;
assign target_only_stripe[2372] = 24'h000000;
assign target_only_stripe[2373] = 24'h000000;
assign target_only_stripe[2374] = 24'h000000;
assign target_only_stripe[2375] = 24'h000000;
assign target_only_stripe[2376] = 24'h000000;
assign target_only_stripe[2377] = 24'h000000;
assign target_only_stripe[2378] = 24'h000000;
assign target_only_stripe[2379] = 24'h000000;
assign target_only_stripe[2380] = 24'h000000;
assign target_only_stripe[2381] = 24'h000000;
assign target_only_stripe[2382] = 24'h000000;
assign target_only_stripe[2383] = 24'h000000;
assign target_only_stripe[2384] = 24'h000000;
assign target_only_stripe[2385] = 24'h000000;
assign target_only_stripe[2386] = 24'h000000;
assign target_only_stripe[2387] = 24'h000000;
assign target_only_stripe[2388] = 24'h000000;
assign target_only_stripe[2389] = 24'h000000;
assign target_only_stripe[2390] = 24'h000000;
assign target_only_stripe[2391] = 24'h000000;
assign target_only_stripe[2392] = 24'h000000;
assign target_only_stripe[2393] = 24'h000000;
assign target_only_stripe[2394] = 24'h000000;
assign target_only_stripe[2395] = 24'h000000;
assign target_only_stripe[2396] = 24'h000000;
assign target_only_stripe[2397] = 24'h000000;
assign target_only_stripe[2398] = 24'h000000;
assign target_only_stripe[2399] = 24'h000000;
assign target_only_stripe[2400] = 24'h000000;
assign target_only_stripe[2401] = 24'h9f9f9f;
assign target_only_stripe[2402] = 24'hffffff;
assign target_only_stripe[2403] = 24'hffffff;
assign target_only_stripe[2404] = 24'hffffff;
assign target_only_stripe[2405] = 24'hffffff;
assign target_only_stripe[2406] = 24'hffffff;
assign target_only_stripe[2407] = 24'hffffff;
assign target_only_stripe[2408] = 24'hffffff;
assign target_only_stripe[2409] = 24'hffffff;
assign target_only_stripe[2410] = 24'hffffff;
assign target_only_stripe[2411] = 24'hffffff;
assign target_only_stripe[2412] = 24'hffffff;
assign target_only_stripe[2413] = 24'hffffff;
assign target_only_stripe[2414] = 24'hffffff;
assign target_only_stripe[2415] = 24'hffffff;
assign target_only_stripe[2416] = 24'hffffff;
assign target_only_stripe[2417] = 24'hffffff;
assign target_only_stripe[2418] = 24'hffffff;
assign target_only_stripe[2419] = 24'hffffff;
assign target_only_stripe[2420] = 24'hffffff;
assign target_only_stripe[2421] = 24'hffffff;
assign target_only_stripe[2422] = 24'hffffff;
assign target_only_stripe[2423] = 24'hffffff;
assign target_only_stripe[2424] = 24'hffffff;
assign target_only_stripe[2425] = 24'hffffff;
assign target_only_stripe[2426] = 24'hffffff;
assign target_only_stripe[2427] = 24'hffffff;
assign target_only_stripe[2428] = 24'hffffff;
assign target_only_stripe[2429] = 24'hffffff;
assign target_only_stripe[2430] = 24'hffffff;
assign target_only_stripe[2431] = 24'hffffff;
assign target_only_stripe[2432] = 24'hffffff;
assign target_only_stripe[2433] = 24'hffffff;
assign target_only_stripe[2434] = 24'hffffff;
assign target_only_stripe[2435] = 24'hffffff;
assign target_only_stripe[2436] = 24'h000000;
assign target_only_stripe[2437] = 24'h000000;
assign target_only_stripe[2438] = 24'h000000;
assign target_only_stripe[2439] = 24'h000000;
assign target_only_stripe[2440] = 24'h000000;
assign target_only_stripe[2441] = 24'h000000;
assign target_only_stripe[2442] = 24'h000000;
assign target_only_stripe[2443] = 24'h000000;
assign target_only_stripe[2444] = 24'h000000;
assign target_only_stripe[2445] = 24'h000000;
assign target_only_stripe[2446] = 24'h000000;
assign target_only_stripe[2447] = 24'h000000;
assign target_only_stripe[2448] = 24'h000000;
assign target_only_stripe[2449] = 24'h000000;
assign target_only_stripe[2450] = 24'h000000;
assign target_only_stripe[2451] = 24'h000000;
assign target_only_stripe[2452] = 24'h000000;
assign target_only_stripe[2453] = 24'h000000;
assign target_only_stripe[2454] = 24'h000000;
assign target_only_stripe[2455] = 24'h000000;
assign target_only_stripe[2456] = 24'h000000;
assign target_only_stripe[2457] = 24'h000000;
assign target_only_stripe[2458] = 24'h000000;
assign target_only_stripe[2459] = 24'h000000;
assign target_only_stripe[2460] = 24'h000000;
assign target_only_stripe[2461] = 24'h000000;
assign target_only_stripe[2462] = 24'h000000;
assign target_only_stripe[2463] = 24'h000000;
assign target_only_stripe[2464] = 24'h000000;
assign target_only_stripe[2465] = 24'h000000;
assign target_only_stripe[2466] = 24'h000000;
assign target_only_stripe[2467] = 24'h000000;
assign target_only_stripe[2468] = 24'h000000;
assign target_only_stripe[2469] = 24'h000000;
assign target_only_stripe[2470] = 24'h000000;
assign target_only_stripe[2471] = 24'h000000;
assign target_only_stripe[2472] = 24'h000000;
assign target_only_stripe[2473] = 24'h000000;
assign target_only_stripe[2474] = 24'h000000;
assign target_only_stripe[2475] = 24'h000000;
assign target_only_stripe[2476] = 24'h000000;
assign target_only_stripe[2477] = 24'h000000;
assign target_only_stripe[2478] = 24'h000000;
assign target_only_stripe[2479] = 24'h000000;
assign target_only_stripe[2480] = 24'h000000;
assign target_only_stripe[2481] = 24'h000000;
assign target_only_stripe[2482] = 24'h000000;
assign target_only_stripe[2483] = 24'h000000;
assign target_only_stripe[2484] = 24'h000000;
assign target_only_stripe[2485] = 24'h000000;
assign target_only_stripe[2486] = 24'h000000;
assign target_only_stripe[2487] = 24'h000000;
assign target_only_stripe[2488] = 24'h000000;
assign target_only_stripe[2489] = 24'h000000;
assign target_only_stripe[2490] = 24'h000000;
assign target_only_stripe[2491] = 24'h000000;
assign target_only_stripe[2492] = 24'h000000;
assign target_only_stripe[2493] = 24'h000000;
assign target_only_stripe[2494] = 24'h000000;
assign target_only_stripe[2495] = 24'h000000;
assign target_only_stripe[2496] = 24'h000000;
assign target_only_stripe[2497] = 24'h000000;
assign target_only_stripe[2498] = 24'h000000;
assign target_only_stripe[2499] = 24'hffffff;
assign target_only_stripe[2500] = 24'hffffff;
assign target_only_stripe[2501] = 24'hffffff;
assign target_only_stripe[2502] = 24'hffffff;
assign target_only_stripe[2503] = 24'hffffff;
assign target_only_stripe[2504] = 24'hffffff;
assign target_only_stripe[2505] = 24'hffffff;
assign target_only_stripe[2506] = 24'hffffff;
assign target_only_stripe[2507] = 24'hffffff;
assign target_only_stripe[2508] = 24'hffffff;
assign target_only_stripe[2509] = 24'hffffff;
assign target_only_stripe[2510] = 24'hffffff;
assign target_only_stripe[2511] = 24'hffffff;
assign target_only_stripe[2512] = 24'hffffff;
assign target_only_stripe[2513] = 24'hffffff;
assign target_only_stripe[2514] = 24'hffffff;
assign target_only_stripe[2515] = 24'hffffff;
assign target_only_stripe[2516] = 24'hffffff;
assign target_only_stripe[2517] = 24'hffffff;
assign target_only_stripe[2518] = 24'hffffff;
assign target_only_stripe[2519] = 24'hffffff;
assign target_only_stripe[2520] = 24'hffffff;
assign target_only_stripe[2521] = 24'hffffff;
assign target_only_stripe[2522] = 24'hffffff;
assign target_only_stripe[2523] = 24'hffffff;
assign target_only_stripe[2524] = 24'hffffff;
assign target_only_stripe[2525] = 24'hffffff;
assign target_only_stripe[2526] = 24'hffffff;
assign target_only_stripe[2527] = 24'hffffff;
assign target_only_stripe[2528] = 24'hffffff;
assign target_only_stripe[2529] = 24'hffffff;
assign target_only_stripe[2530] = 24'hffffff;
assign target_only_stripe[2531] = 24'hffffff;
assign target_only_stripe[2532] = 24'hffffff;
assign target_only_stripe[2533] = 24'h909090;
assign target_only_stripe[2534] = 24'h000000;
assign target_only_stripe[2535] = 24'h000000;
assign target_only_stripe[2536] = 24'h000000;
assign target_only_stripe[2537] = 24'h000000;
assign target_only_stripe[2538] = 24'h000000;
assign target_only_stripe[2539] = 24'h000000;
assign target_only_stripe[2540] = 24'h000000;
assign target_only_stripe[2541] = 24'h000000;
assign target_only_stripe[2542] = 24'h000000;
assign target_only_stripe[2543] = 24'h000000;
assign target_only_stripe[2544] = 24'h000000;
assign target_only_stripe[2545] = 24'h000000;
assign target_only_stripe[2546] = 24'h000000;
assign target_only_stripe[2547] = 24'h000000;
assign target_only_stripe[2548] = 24'h000000;
assign target_only_stripe[2549] = 24'h000000;
assign target_only_stripe[2550] = 24'h000000;
assign target_only_stripe[2551] = 24'h000000;
assign target_only_stripe[2552] = 24'h000000;
assign target_only_stripe[2553] = 24'h000000;
assign target_only_stripe[2554] = 24'h000000;
assign target_only_stripe[2555] = 24'h000000;
assign target_only_stripe[2556] = 24'h000000;
assign target_only_stripe[2557] = 24'h000000;
assign target_only_stripe[2558] = 24'h000000;
assign target_only_stripe[2559] = 24'h000000;
assign target_only_stripe[2560] = 24'h000000;
assign target_only_stripe[2561] = 24'h000000;
assign target_only_stripe[2562] = 24'h000000;
assign target_only_stripe[2563] = 24'h000000;
assign target_only_stripe[2564] = 24'h000000;
assign target_only_stripe[2565] = 24'h000000;
assign target_only_stripe[2566] = 24'hb7b7b7;
assign target_only_stripe[2567] = 24'hffffff;
assign target_only_stripe[2568] = 24'hffffff;
assign target_only_stripe[2569] = 24'hffffff;
assign target_only_stripe[2570] = 24'hffffff;
assign target_only_stripe[2571] = 24'hffffff;
assign target_only_stripe[2572] = 24'hffffff;
assign target_only_stripe[2573] = 24'hffffff;
assign target_only_stripe[2574] = 24'hffffff;
assign target_only_stripe[2575] = 24'hffffff;
assign target_only_stripe[2576] = 24'hffffff;
assign target_only_stripe[2577] = 24'hffffff;
assign target_only_stripe[2578] = 24'hffffff;
assign target_only_stripe[2579] = 24'hffffff;
assign target_only_stripe[2580] = 24'hffffff;
assign target_only_stripe[2581] = 24'hffffff;
assign target_only_stripe[2582] = 24'hffffff;
assign target_only_stripe[2583] = 24'hffffff;
assign target_only_stripe[2584] = 24'hffffff;
assign target_only_stripe[2585] = 24'hffffff;
assign target_only_stripe[2586] = 24'hffffff;
assign target_only_stripe[2587] = 24'hffffff;
assign target_only_stripe[2588] = 24'hffffff;
assign target_only_stripe[2589] = 24'hffffff;
assign target_only_stripe[2590] = 24'hffffff;
assign target_only_stripe[2591] = 24'hffffff;
assign target_only_stripe[2592] = 24'hffffff;
assign target_only_stripe[2593] = 24'hffffff;
assign target_only_stripe[2594] = 24'hffffff;
assign target_only_stripe[2595] = 24'hffffff;
assign target_only_stripe[2596] = 24'hffffff;
assign target_only_stripe[2597] = 24'hffffff;
assign target_only_stripe[2598] = 24'hffffff;
assign target_only_stripe[2599] = 24'he1d8d5;
assign target_only_stripe[2600] = 24'h1b1b1b;
assign target_only_stripe[2601] = 24'h000000;
assign target_only_stripe[2602] = 24'h000000;
assign target_only_stripe[2603] = 24'h000000;
assign target_only_stripe[2604] = 24'h000000;
assign target_only_stripe[2605] = 24'h000000;
assign target_only_stripe[2606] = 24'h000000;
assign target_only_stripe[2607] = 24'h000000;
assign target_only_stripe[2608] = 24'h000000;
assign target_only_stripe[2609] = 24'h000000;
assign target_only_stripe[2610] = 24'h000000;
assign target_only_stripe[2611] = 24'h000000;
assign target_only_stripe[2612] = 24'h000000;
assign target_only_stripe[2613] = 24'h000000;
assign target_only_stripe[2614] = 24'h000000;
assign target_only_stripe[2615] = 24'h000000;
assign target_only_stripe[2616] = 24'h000000;
assign target_only_stripe[2617] = 24'h000000;
assign target_only_stripe[2618] = 24'h000000;
assign target_only_stripe[2619] = 24'h000000;
assign target_only_stripe[2620] = 24'h000000;
assign target_only_stripe[2621] = 24'h000000;
assign target_only_stripe[2622] = 24'h000000;
assign target_only_stripe[2623] = 24'h000000;
assign target_only_stripe[2624] = 24'h000000;
assign target_only_stripe[2625] = 24'h000000;
assign target_only_stripe[2626] = 24'h000000;
assign target_only_stripe[2627] = 24'h000000;
assign target_only_stripe[2628] = 24'h000000;
assign target_only_stripe[2629] = 24'h000000;
assign target_only_stripe[2630] = 24'h000000;
assign target_only_stripe[2631] = 24'h000000;
assign target_only_stripe[2632] = 24'h000000;
assign target_only_stripe[2633] = 24'h000000;
assign target_only_stripe[2634] = 24'h000000;
assign target_only_stripe[2635] = 24'h000000;
assign target_only_stripe[2636] = 24'h000000;
assign target_only_stripe[2637] = 24'h000000;
assign target_only_stripe[2638] = 24'h000000;
assign target_only_stripe[2639] = 24'h000000;
assign target_only_stripe[2640] = 24'h000000;
assign target_only_stripe[2641] = 24'h000000;
assign target_only_stripe[2642] = 24'h000000;
assign target_only_stripe[2643] = 24'h000000;
assign target_only_stripe[2644] = 24'h000000;
assign target_only_stripe[2645] = 24'h000000;
assign target_only_stripe[2646] = 24'h000000;
assign target_only_stripe[2647] = 24'h000000;
assign target_only_stripe[2648] = 24'h000000;
assign target_only_stripe[2649] = 24'h000000;
assign target_only_stripe[2650] = 24'h000000;
assign target_only_stripe[2651] = 24'h000000;
assign target_only_stripe[2652] = 24'h000000;
assign target_only_stripe[2653] = 24'h000000;
assign target_only_stripe[2654] = 24'h000000;
assign target_only_stripe[2655] = 24'h000000;
assign target_only_stripe[2656] = 24'h000000;
assign target_only_stripe[2657] = 24'h000000;
assign target_only_stripe[2658] = 24'h000000;
assign target_only_stripe[2659] = 24'h000000;
assign target_only_stripe[2660] = 24'h000000;
assign target_only_stripe[2661] = 24'h000000;
assign target_only_stripe[2662] = 24'h000000;
assign target_only_stripe[2663] = 24'h121212;
assign target_only_stripe[2664] = 24'he9e7e6;
assign target_only_stripe[2665] = 24'hffffff;
assign target_only_stripe[2666] = 24'hffffff;
assign target_only_stripe[2667] = 24'hffffff;
assign target_only_stripe[2668] = 24'hffffff;
assign target_only_stripe[2669] = 24'hffffff;
assign target_only_stripe[2670] = 24'hffffff;
assign target_only_stripe[2671] = 24'hffffff;
assign target_only_stripe[2672] = 24'hffffff;
assign target_only_stripe[2673] = 24'hffffff;
assign target_only_stripe[2674] = 24'hffffff;
assign target_only_stripe[2675] = 24'hffffff;
assign target_only_stripe[2676] = 24'hffffff;
assign target_only_stripe[2677] = 24'hffffff;
assign target_only_stripe[2678] = 24'hffffff;
assign target_only_stripe[2679] = 24'hffffff;
assign target_only_stripe[2680] = 24'hffffff;
assign target_only_stripe[2681] = 24'hffffff;
assign target_only_stripe[2682] = 24'hffffff;
assign target_only_stripe[2683] = 24'hffffff;
assign target_only_stripe[2684] = 24'hffffff;
assign target_only_stripe[2685] = 24'hffffff;
assign target_only_stripe[2686] = 24'hffffff;
assign target_only_stripe[2687] = 24'hffffff;
assign target_only_stripe[2688] = 24'hffffff;
assign target_only_stripe[2689] = 24'hffffff;
assign target_only_stripe[2690] = 24'hffffff;
assign target_only_stripe[2691] = 24'hffffff;
assign target_only_stripe[2692] = 24'hffffff;
assign target_only_stripe[2693] = 24'hffffff;
assign target_only_stripe[2694] = 24'hfaf7f5;
assign target_only_stripe[2695] = 24'hffffff;
assign target_only_stripe[2696] = 24'hffffff;
assign target_only_stripe[2697] = 24'haaaaaa;
assign target_only_stripe[2698] = 24'h000000;
assign target_only_stripe[2699] = 24'h000000;
assign target_only_stripe[2700] = 24'h000000;
assign target_only_stripe[2701] = 24'h000000;
assign target_only_stripe[2702] = 24'h000000;
assign target_only_stripe[2703] = 24'h000000;
assign target_only_stripe[2704] = 24'h000000;
assign target_only_stripe[2705] = 24'h000000;
assign target_only_stripe[2706] = 24'h000000;
assign target_only_stripe[2707] = 24'h000000;
assign target_only_stripe[2708] = 24'h000000;
assign target_only_stripe[2709] = 24'h000000;
assign target_only_stripe[2710] = 24'h000000;
assign target_only_stripe[2711] = 24'h000000;
assign target_only_stripe[2712] = 24'h000000;
assign target_only_stripe[2713] = 24'h000000;
assign target_only_stripe[2714] = 24'h000000;
assign target_only_stripe[2715] = 24'h000000;
assign target_only_stripe[2716] = 24'h000000;
assign target_only_stripe[2717] = 24'h000000;
assign target_only_stripe[2718] = 24'h000000;
assign target_only_stripe[2719] = 24'h000000;
assign target_only_stripe[2720] = 24'h000000;
assign target_only_stripe[2721] = 24'h000000;
assign target_only_stripe[2722] = 24'h000000;
assign target_only_stripe[2723] = 24'h000000;
assign target_only_stripe[2724] = 24'h000000;
assign target_only_stripe[2725] = 24'h000000;
assign target_only_stripe[2726] = 24'h000000;
assign target_only_stripe[2727] = 24'h000000;
assign target_only_stripe[2728] = 24'h000000;
assign target_only_stripe[2729] = 24'h000000;
assign target_only_stripe[2730] = 24'h949494;
assign target_only_stripe[2731] = 24'hffffff;
assign target_only_stripe[2732] = 24'hffffff;
assign target_only_stripe[2733] = 24'hffffff;
assign target_only_stripe[2734] = 24'hffffff;
assign target_only_stripe[2735] = 24'hffffff;
assign target_only_stripe[2736] = 24'hffffff;
assign target_only_stripe[2737] = 24'hffffff;
assign target_only_stripe[2738] = 24'hffffff;
assign target_only_stripe[2739] = 24'hffffff;
assign target_only_stripe[2740] = 24'hffffff;
assign target_only_stripe[2741] = 24'hffffff;
assign target_only_stripe[2742] = 24'hffffff;
assign target_only_stripe[2743] = 24'hffffff;
assign target_only_stripe[2744] = 24'hffffff;
assign target_only_stripe[2745] = 24'hffffff;
assign target_only_stripe[2746] = 24'hffffff;
assign target_only_stripe[2747] = 24'hffffff;
assign target_only_stripe[2748] = 24'hffffff;
assign target_only_stripe[2749] = 24'hffffff;
assign target_only_stripe[2750] = 24'hffffff;
assign target_only_stripe[2751] = 24'hffffff;
assign target_only_stripe[2752] = 24'hffffff;
assign target_only_stripe[2753] = 24'hffffff;
assign target_only_stripe[2754] = 24'hffffff;
assign target_only_stripe[2755] = 24'hffffff;
assign target_only_stripe[2756] = 24'hffffff;
assign target_only_stripe[2757] = 24'hffffff;
assign target_only_stripe[2758] = 24'hffffff;
assign target_only_stripe[2759] = 24'hffffff;
assign target_only_stripe[2760] = 24'hffffff;
assign target_only_stripe[2761] = 24'hffffff;
assign target_only_stripe[2762] = 24'hffffff;
assign target_only_stripe[2763] = 24'hffffff;
assign target_only_stripe[2764] = 24'hffffff;
assign target_only_stripe[2765] = 24'h000000;
assign target_only_stripe[2766] = 24'h000000;
assign target_only_stripe[2767] = 24'h000000;
assign target_only_stripe[2768] = 24'h000000;
assign target_only_stripe[2769] = 24'h000000;
assign target_only_stripe[2770] = 24'h000000;
assign target_only_stripe[2771] = 24'h000000;
assign target_only_stripe[2772] = 24'h000000;
assign target_only_stripe[2773] = 24'h000000;
assign target_only_stripe[2774] = 24'h000000;
assign target_only_stripe[2775] = 24'h000000;
assign target_only_stripe[2776] = 24'h000000;
assign target_only_stripe[2777] = 24'h000000;
assign target_only_stripe[2778] = 24'h000000;
assign target_only_stripe[2779] = 24'h000000;
assign target_only_stripe[2780] = 24'h000000;
assign target_only_stripe[2781] = 24'h000000;
assign target_only_stripe[2782] = 24'h000000;
assign target_only_stripe[2783] = 24'h000000;
assign target_only_stripe[2784] = 24'h000000;
assign target_only_stripe[2785] = 24'h000000;
assign target_only_stripe[2786] = 24'h000000;
assign target_only_stripe[2787] = 24'h000000;
assign target_only_stripe[2788] = 24'h000000;
assign target_only_stripe[2789] = 24'h000000;
assign target_only_stripe[2790] = 24'h000000;
assign target_only_stripe[2791] = 24'h000000;
assign target_only_stripe[2792] = 24'h000000;
assign target_only_stripe[2793] = 24'h000000;
assign target_only_stripe[2794] = 24'h000000;
assign target_only_stripe[2795] = 24'h000000;
assign target_only_stripe[2796] = 24'h000000;
assign target_only_stripe[2797] = 24'h000000;
assign target_only_stripe[2798] = 24'h000000;
assign target_only_stripe[2799] = 24'h000000;
assign target_only_stripe[2800] = 24'h000000;
assign target_only_stripe[2801] = 24'h000000;
assign target_only_stripe[2802] = 24'h000000;
assign target_only_stripe[2803] = 24'h000000;
assign target_only_stripe[2804] = 24'h000000;
assign target_only_stripe[2805] = 24'h000000;
assign target_only_stripe[2806] = 24'h000000;
assign target_only_stripe[2807] = 24'h000000;
assign target_only_stripe[2808] = 24'h000000;
assign target_only_stripe[2809] = 24'h000000;
assign target_only_stripe[2810] = 24'h000000;
assign target_only_stripe[2811] = 24'h000000;
assign target_only_stripe[2812] = 24'h000000;
assign target_only_stripe[2813] = 24'h000000;
assign target_only_stripe[2814] = 24'h000000;
assign target_only_stripe[2815] = 24'h000000;
assign target_only_stripe[2816] = 24'h000000;
assign target_only_stripe[2817] = 24'h000000;
assign target_only_stripe[2818] = 24'h000000;
assign target_only_stripe[2819] = 24'h000000;
assign target_only_stripe[2820] = 24'h000000;
assign target_only_stripe[2821] = 24'h000000;
assign target_only_stripe[2822] = 24'h000000;
assign target_only_stripe[2823] = 24'h000000;
assign target_only_stripe[2824] = 24'h000000;
assign target_only_stripe[2825] = 24'h000000;
assign target_only_stripe[2826] = 24'h000000;
assign target_only_stripe[2827] = 24'h000000;
assign target_only_stripe[2828] = 24'hffffff;
assign target_only_stripe[2829] = 24'hffffff;
assign target_only_stripe[2830] = 24'hffffff;
assign target_only_stripe[2831] = 24'hffffff;
assign target_only_stripe[2832] = 24'hffffff;
assign target_only_stripe[2833] = 24'hffffff;
assign target_only_stripe[2834] = 24'hffffff;
assign target_only_stripe[2835] = 24'hffffff;
assign target_only_stripe[2836] = 24'hffffff;
assign target_only_stripe[2837] = 24'hffffff;
assign target_only_stripe[2838] = 24'hffffff;
assign target_only_stripe[2839] = 24'hffffff;
assign target_only_stripe[2840] = 24'hffffff;
assign target_only_stripe[2841] = 24'hffffff;
assign target_only_stripe[2842] = 24'hffffff;
assign target_only_stripe[2843] = 24'hffffff;
assign target_only_stripe[2844] = 24'hffffff;
assign target_only_stripe[2845] = 24'hffffff;
assign target_only_stripe[2846] = 24'hffffff;
assign target_only_stripe[2847] = 24'hffffff;
assign target_only_stripe[2848] = 24'hffffff;
assign target_only_stripe[2849] = 24'hffffff;
assign target_only_stripe[2850] = 24'hffffff;
assign target_only_stripe[2851] = 24'hffffff;
assign target_only_stripe[2852] = 24'hffffff;
assign target_only_stripe[2853] = 24'hffffff;
assign target_only_stripe[2854] = 24'hffffff;
assign target_only_stripe[2855] = 24'hffffff;
assign target_only_stripe[2856] = 24'hffffff;
assign target_only_stripe[2857] = 24'hffffff;
assign target_only_stripe[2858] = 24'hffffff;
assign target_only_stripe[2859] = 24'hffffff;
assign target_only_stripe[2860] = 24'hffffff;
assign target_only_stripe[2861] = 24'hffffff;
assign target_only_stripe[2862] = 24'h9c9c9c;
assign target_only_stripe[2863] = 24'h000000;
assign target_only_stripe[2864] = 24'h000000;
assign target_only_stripe[2865] = 24'h000000;
assign target_only_stripe[2866] = 24'h000000;
assign target_only_stripe[2867] = 24'h000000;
assign target_only_stripe[2868] = 24'h000000;
assign target_only_stripe[2869] = 24'h000000;
assign target_only_stripe[2870] = 24'h000000;
assign target_only_stripe[2871] = 24'h000000;
assign target_only_stripe[2872] = 24'h000000;
assign target_only_stripe[2873] = 24'h000000;
assign target_only_stripe[2874] = 24'h000000;
assign target_only_stripe[2875] = 24'h000000;
assign target_only_stripe[2876] = 24'h000000;
assign target_only_stripe[2877] = 24'h000000;
assign target_only_stripe[2878] = 24'h000000;
assign target_only_stripe[2879] = 24'h000000;
assign target_only_stripe[2880] = 24'h000000;
assign target_only_stripe[2881] = 24'h000000;
assign target_only_stripe[2882] = 24'h000000;
assign target_only_stripe[2883] = 24'h000000;
assign target_only_stripe[2884] = 24'h000000;
assign target_only_stripe[2885] = 24'h000000;
assign target_only_stripe[2886] = 24'h000000;
assign target_only_stripe[2887] = 24'h000000;
assign target_only_stripe[2888] = 24'h000000;
assign target_only_stripe[2889] = 24'h000000;
assign target_only_stripe[2890] = 24'h000000;
assign target_only_stripe[2891] = 24'h000000;
assign target_only_stripe[2892] = 24'h000000;
assign target_only_stripe[2893] = 24'h000000;
assign target_only_stripe[2894] = 24'h000000;
assign target_only_stripe[2895] = 24'ha3a3a3;
assign target_only_stripe[2896] = 24'hffffff;
assign target_only_stripe[2897] = 24'hffffff;
assign target_only_stripe[2898] = 24'hffffff;
assign target_only_stripe[2899] = 24'hffffff;
assign target_only_stripe[2900] = 24'hffffff;
assign target_only_stripe[2901] = 24'hffffff;
assign target_only_stripe[2902] = 24'hffffff;
assign target_only_stripe[2903] = 24'hffffff;
assign target_only_stripe[2904] = 24'hffffff;
assign target_only_stripe[2905] = 24'hffffff;
assign target_only_stripe[2906] = 24'hffffff;
assign target_only_stripe[2907] = 24'hffffff;
assign target_only_stripe[2908] = 24'hffffff;
assign target_only_stripe[2909] = 24'hffffff;
assign target_only_stripe[2910] = 24'hffffff;
assign target_only_stripe[2911] = 24'hffffff;
assign target_only_stripe[2912] = 24'hffffff;
assign target_only_stripe[2913] = 24'hffffff;
assign target_only_stripe[2914] = 24'hffffff;
assign target_only_stripe[2915] = 24'hffffff;
assign target_only_stripe[2916] = 24'hffffff;
assign target_only_stripe[2917] = 24'hffffff;
assign target_only_stripe[2918] = 24'hffffff;
assign target_only_stripe[2919] = 24'hffffff;
assign target_only_stripe[2920] = 24'hffffff;
assign target_only_stripe[2921] = 24'hffffff;
assign target_only_stripe[2922] = 24'hffffff;
assign target_only_stripe[2923] = 24'hffffff;
assign target_only_stripe[2924] = 24'hffffff;
assign target_only_stripe[2925] = 24'hffffff;
assign target_only_stripe[2926] = 24'hffffff;
assign target_only_stripe[2927] = 24'hffffff;
assign target_only_stripe[2928] = 24'hceb7ab;
assign target_only_stripe[2929] = 24'h1b1b1b;
assign target_only_stripe[2930] = 24'h000000;
assign target_only_stripe[2931] = 24'h000000;
assign target_only_stripe[2932] = 24'h000000;
assign target_only_stripe[2933] = 24'h000000;
assign target_only_stripe[2934] = 24'h000000;
assign target_only_stripe[2935] = 24'h000000;
assign target_only_stripe[2936] = 24'h000000;
assign target_only_stripe[2937] = 24'h000000;
assign target_only_stripe[2938] = 24'h000000;
assign target_only_stripe[2939] = 24'h000000;
assign target_only_stripe[2940] = 24'h000000;
assign target_only_stripe[2941] = 24'h000000;
assign target_only_stripe[2942] = 24'h000000;
assign target_only_stripe[2943] = 24'h000000;
assign target_only_stripe[2944] = 24'h000000;
assign target_only_stripe[2945] = 24'h000000;
assign target_only_stripe[2946] = 24'h000000;
assign target_only_stripe[2947] = 24'h000000;
assign target_only_stripe[2948] = 24'h000000;
assign target_only_stripe[2949] = 24'h000000;
assign target_only_stripe[2950] = 24'h000000;
assign target_only_stripe[2951] = 24'h000000;
assign target_only_stripe[2952] = 24'h000000;
assign target_only_stripe[2953] = 24'h000000;
assign target_only_stripe[2954] = 24'h000000;
assign target_only_stripe[2955] = 24'h000000;
assign target_only_stripe[2956] = 24'h000000;
assign target_only_stripe[2957] = 24'h000000;
assign target_only_stripe[2958] = 24'h000000;
assign target_only_stripe[2959] = 24'h000000;
assign target_only_stripe[2960] = 24'h000000;
assign target_only_stripe[2961] = 24'h000000;
assign target_only_stripe[2962] = 24'h000000;
assign target_only_stripe[2963] = 24'h000000;
assign target_only_stripe[2964] = 24'h000000;
assign target_only_stripe[2965] = 24'h000000;
assign target_only_stripe[2966] = 24'h000000;
assign target_only_stripe[2967] = 24'h000000;
assign target_only_stripe[2968] = 24'h000000;
assign target_only_stripe[2969] = 24'h000000;
assign target_only_stripe[2970] = 24'h000000;
assign target_only_stripe[2971] = 24'h000000;
assign target_only_stripe[2972] = 24'h000000;
assign target_only_stripe[2973] = 24'h000000;
assign target_only_stripe[2974] = 24'h000000;
assign target_only_stripe[2975] = 24'h000000;
assign target_only_stripe[2976] = 24'h000000;
assign target_only_stripe[2977] = 24'h000000;
assign target_only_stripe[2978] = 24'h000000;
assign target_only_stripe[2979] = 24'h000000;
assign target_only_stripe[2980] = 24'h000000;
assign target_only_stripe[2981] = 24'h000000;
assign target_only_stripe[2982] = 24'h000000;
assign target_only_stripe[2983] = 24'h000000;
assign target_only_stripe[2984] = 24'h000000;
assign target_only_stripe[2985] = 24'h000000;
assign target_only_stripe[2986] = 24'h000000;
assign target_only_stripe[2987] = 24'h000000;
assign target_only_stripe[2988] = 24'h000000;
assign target_only_stripe[2989] = 24'h000000;
assign target_only_stripe[2990] = 24'h000000;
assign target_only_stripe[2991] = 24'h000000;
assign target_only_stripe[2992] = 24'h121212;
assign target_only_stripe[2993] = 24'he8e7e6;
assign target_only_stripe[2994] = 24'hffffff;
assign target_only_stripe[2995] = 24'hffffff;
assign target_only_stripe[2996] = 24'hffffff;
assign target_only_stripe[2997] = 24'hffffff;
assign target_only_stripe[2998] = 24'hffffff;
assign target_only_stripe[2999] = 24'hffffff;
assign target_only_stripe[3000] = 24'hffffff;
assign target_only_stripe[3001] = 24'hffffff;
assign target_only_stripe[3002] = 24'hffffff;
assign target_only_stripe[3003] = 24'hffffff;
assign target_only_stripe[3004] = 24'hffffff;
assign target_only_stripe[3005] = 24'hffffff;
assign target_only_stripe[3006] = 24'hffffff;
assign target_only_stripe[3007] = 24'hffffff;
assign target_only_stripe[3008] = 24'hffffff;
assign target_only_stripe[3009] = 24'hffffff;
assign target_only_stripe[3010] = 24'hffffff;
assign target_only_stripe[3011] = 24'hffffff;
assign target_only_stripe[3012] = 24'hffffff;
assign target_only_stripe[3013] = 24'hffffff;
assign target_only_stripe[3014] = 24'hffffff;
assign target_only_stripe[3015] = 24'hffffff;
assign target_only_stripe[3016] = 24'hffffff;
assign target_only_stripe[3017] = 24'hffffff;
assign target_only_stripe[3018] = 24'hffffff;
assign target_only_stripe[3019] = 24'hffffff;
assign target_only_stripe[3020] = 24'hffffff;
assign target_only_stripe[3021] = 24'hffffff;
assign target_only_stripe[3022] = 24'hfaf7f5;
assign target_only_stripe[3023] = 24'hffffff;
assign target_only_stripe[3024] = 24'hffffff;
assign target_only_stripe[3025] = 24'hffffff;
assign target_only_stripe[3026] = 24'h9f9f9f;
assign target_only_stripe[3027] = 24'h000000;
assign target_only_stripe[3028] = 24'h000000;
assign target_only_stripe[3029] = 24'h000000;
assign target_only_stripe[3030] = 24'h000000;
assign target_only_stripe[3031] = 24'h000000;
assign target_only_stripe[3032] = 24'h000000;
assign target_only_stripe[3033] = 24'h000000;
assign target_only_stripe[3034] = 24'h000000;
assign target_only_stripe[3035] = 24'h000000;
assign target_only_stripe[3036] = 24'h000000;
assign target_only_stripe[3037] = 24'h000000;
assign target_only_stripe[3038] = 24'h000000;
assign target_only_stripe[3039] = 24'h000000;
assign target_only_stripe[3040] = 24'h000000;
assign target_only_stripe[3041] = 24'h000000;
assign target_only_stripe[3042] = 24'h000000;
assign target_only_stripe[3043] = 24'h000000;
assign target_only_stripe[3044] = 24'h000000;
assign target_only_stripe[3045] = 24'h000000;
assign target_only_stripe[3046] = 24'h000000;
assign target_only_stripe[3047] = 24'h000000;
assign target_only_stripe[3048] = 24'h000000;
assign target_only_stripe[3049] = 24'h000000;
assign target_only_stripe[3050] = 24'h000000;
assign target_only_stripe[3051] = 24'h000000;
assign target_only_stripe[3052] = 24'h000000;
assign target_only_stripe[3053] = 24'h000000;
assign target_only_stripe[3054] = 24'h000000;
assign target_only_stripe[3055] = 24'h000000;
assign target_only_stripe[3056] = 24'h000000;
assign target_only_stripe[3057] = 24'h000000;
assign target_only_stripe[3058] = 24'h000000;
assign target_only_stripe[3059] = 24'h999999;
assign target_only_stripe[3060] = 24'hffffff;
assign target_only_stripe[3061] = 24'hffffff;
assign target_only_stripe[3062] = 24'hffffff;
assign target_only_stripe[3063] = 24'hffffff;
assign target_only_stripe[3064] = 24'hffffff;
assign target_only_stripe[3065] = 24'hffffff;
assign target_only_stripe[3066] = 24'hffffff;
assign target_only_stripe[3067] = 24'hffffff;
assign target_only_stripe[3068] = 24'hffffff;
assign target_only_stripe[3069] = 24'hffffff;
assign target_only_stripe[3070] = 24'hffffff;
assign target_only_stripe[3071] = 24'hffffff;
assign target_only_stripe[3072] = 24'hffffff;
assign target_only_stripe[3073] = 24'hffffff;
assign target_only_stripe[3074] = 24'hffffff;
assign target_only_stripe[3075] = 24'hffffff;
assign target_only_stripe[3076] = 24'hffffff;
assign target_only_stripe[3077] = 24'hffffff;
assign target_only_stripe[3078] = 24'hffffff;
assign target_only_stripe[3079] = 24'hffffff;
assign target_only_stripe[3080] = 24'hffffff;
assign target_only_stripe[3081] = 24'hffffff;
assign target_only_stripe[3082] = 24'hffffff;
assign target_only_stripe[3083] = 24'hffffff;
assign target_only_stripe[3084] = 24'hffffff;
assign target_only_stripe[3085] = 24'hffffff;
assign target_only_stripe[3086] = 24'hffffff;
assign target_only_stripe[3087] = 24'hffffff;
assign target_only_stripe[3088] = 24'hffffff;
assign target_only_stripe[3089] = 24'hffffff;
assign target_only_stripe[3090] = 24'hffffff;
assign target_only_stripe[3091] = 24'hffffff;
assign target_only_stripe[3092] = 24'hffffff;
assign target_only_stripe[3093] = 24'h9e9e9e;
assign target_only_stripe[3094] = 24'h000000;
assign target_only_stripe[3095] = 24'h000000;
assign target_only_stripe[3096] = 24'h000000;
assign target_only_stripe[3097] = 24'h000000;
assign target_only_stripe[3098] = 24'h000000;
assign target_only_stripe[3099] = 24'h000000;
assign target_only_stripe[3100] = 24'h000000;
assign target_only_stripe[3101] = 24'h000000;
assign target_only_stripe[3102] = 24'h000000;
assign target_only_stripe[3103] = 24'h000000;
assign target_only_stripe[3104] = 24'h000000;
assign target_only_stripe[3105] = 24'h000000;
assign target_only_stripe[3106] = 24'h000000;
assign target_only_stripe[3107] = 24'h000000;
assign target_only_stripe[3108] = 24'h000000;
assign target_only_stripe[3109] = 24'h000000;
assign target_only_stripe[3110] = 24'h000000;
assign target_only_stripe[3111] = 24'h000000;
assign target_only_stripe[3112] = 24'h000000;
assign target_only_stripe[3113] = 24'h000000;
assign target_only_stripe[3114] = 24'h000000;
assign target_only_stripe[3115] = 24'h000000;
assign target_only_stripe[3116] = 24'h000000;
assign target_only_stripe[3117] = 24'h000000;
assign target_only_stripe[3118] = 24'h000000;
assign target_only_stripe[3119] = 24'h000000;
assign target_only_stripe[3120] = 24'h000000;
assign target_only_stripe[3121] = 24'h000000;
assign target_only_stripe[3122] = 24'h000000;
assign target_only_stripe[3123] = 24'h000000;
assign target_only_stripe[3124] = 24'h000000;
assign target_only_stripe[3125] = 24'h000000;
assign target_only_stripe[3126] = 24'h000000;
assign target_only_stripe[3127] = 24'h000000;
assign target_only_stripe[3128] = 24'h000000;
assign target_only_stripe[3129] = 24'h000000;
assign target_only_stripe[3130] = 24'h000000;
assign target_only_stripe[3131] = 24'h000000;
assign target_only_stripe[3132] = 24'h000000;
assign target_only_stripe[3133] = 24'h000000;
assign target_only_stripe[3134] = 24'h000000;
assign target_only_stripe[3135] = 24'h000000;
assign target_only_stripe[3136] = 24'h000000;
assign target_only_stripe[3137] = 24'h000000;
assign target_only_stripe[3138] = 24'h000000;
assign target_only_stripe[3139] = 24'h000000;
assign target_only_stripe[3140] = 24'h000000;
assign target_only_stripe[3141] = 24'h000000;
assign target_only_stripe[3142] = 24'h000000;
assign target_only_stripe[3143] = 24'h000000;
assign target_only_stripe[3144] = 24'h000000;
assign target_only_stripe[3145] = 24'h000000;
assign target_only_stripe[3146] = 24'h000000;
assign target_only_stripe[3147] = 24'h000000;
assign target_only_stripe[3148] = 24'h000000;
assign target_only_stripe[3149] = 24'h000000;
assign target_only_stripe[3150] = 24'h000000;
assign target_only_stripe[3151] = 24'h000000;
assign target_only_stripe[3152] = 24'h000000;
assign target_only_stripe[3153] = 24'h000000;
assign target_only_stripe[3154] = 24'h000000;
assign target_only_stripe[3155] = 24'h000000;
assign target_only_stripe[3156] = 24'h000000;
assign target_only_stripe[3157] = 24'h434343;
assign target_only_stripe[3158] = 24'hffffff;
assign target_only_stripe[3159] = 24'hffffff;
assign target_only_stripe[3160] = 24'hffffff;
assign target_only_stripe[3161] = 24'hffffff;
assign target_only_stripe[3162] = 24'hffffff;
assign target_only_stripe[3163] = 24'hffffff;
assign target_only_stripe[3164] = 24'hffffff;
assign target_only_stripe[3165] = 24'hffffff;
assign target_only_stripe[3166] = 24'hffffff;
assign target_only_stripe[3167] = 24'hffffff;
assign target_only_stripe[3168] = 24'hffffff;
assign target_only_stripe[3169] = 24'hffffff;
assign target_only_stripe[3170] = 24'hffffff;
assign target_only_stripe[3171] = 24'hffffff;
assign target_only_stripe[3172] = 24'hffffff;
assign target_only_stripe[3173] = 24'hffffff;
assign target_only_stripe[3174] = 24'hffffff;
assign target_only_stripe[3175] = 24'hffffff;
assign target_only_stripe[3176] = 24'hffffff;
assign target_only_stripe[3177] = 24'hffffff;
assign target_only_stripe[3178] = 24'hffffff;
assign target_only_stripe[3179] = 24'hffffff;
assign target_only_stripe[3180] = 24'hffffff;
assign target_only_stripe[3181] = 24'hffffff;
assign target_only_stripe[3182] = 24'hffffff;
assign target_only_stripe[3183] = 24'hffffff;
assign target_only_stripe[3184] = 24'hffffff;
assign target_only_stripe[3185] = 24'hffffff;
assign target_only_stripe[3186] = 24'hffffff;
assign target_only_stripe[3187] = 24'hffffff;
assign target_only_stripe[3188] = 24'hffffff;
assign target_only_stripe[3189] = 24'hffffff;
assign target_only_stripe[3190] = 24'hffffff;
assign target_only_stripe[3191] = 24'ha1a1a1;
assign target_only_stripe[3192] = 24'h000000;
assign target_only_stripe[3193] = 24'h000000;
assign target_only_stripe[3194] = 24'h000000;
assign target_only_stripe[3195] = 24'h000000;
assign target_only_stripe[3196] = 24'h000000;
assign target_only_stripe[3197] = 24'h000000;
assign target_only_stripe[3198] = 24'h000000;
assign target_only_stripe[3199] = 24'h000000;
assign target_only_stripe[3200] = 24'h000000;
assign target_only_stripe[3201] = 24'h000000;
assign target_only_stripe[3202] = 24'h000000;
assign target_only_stripe[3203] = 24'h000000;
assign target_only_stripe[3204] = 24'h000000;
assign target_only_stripe[3205] = 24'h000000;
assign target_only_stripe[3206] = 24'h000000;
assign target_only_stripe[3207] = 24'h000000;
assign target_only_stripe[3208] = 24'h000000;
assign target_only_stripe[3209] = 24'h000000;
assign target_only_stripe[3210] = 24'h000000;
assign target_only_stripe[3211] = 24'h000000;
assign target_only_stripe[3212] = 24'h000000;
assign target_only_stripe[3213] = 24'h000000;
assign target_only_stripe[3214] = 24'h000000;
assign target_only_stripe[3215] = 24'h000000;
assign target_only_stripe[3216] = 24'h000000;
assign target_only_stripe[3217] = 24'h000000;
assign target_only_stripe[3218] = 24'h000000;
assign target_only_stripe[3219] = 24'h000000;
assign target_only_stripe[3220] = 24'h000000;
assign target_only_stripe[3221] = 24'h000000;
assign target_only_stripe[3222] = 24'h000000;
assign target_only_stripe[3223] = 24'h000000;
assign target_only_stripe[3224] = 24'hb5b5b5;
assign target_only_stripe[3225] = 24'hffffff;
assign target_only_stripe[3226] = 24'hffffff;
assign target_only_stripe[3227] = 24'hffffff;
assign target_only_stripe[3228] = 24'hffffff;
assign target_only_stripe[3229] = 24'hffffff;
assign target_only_stripe[3230] = 24'hffffff;
assign target_only_stripe[3231] = 24'hffffff;
assign target_only_stripe[3232] = 24'hffffff;
assign target_only_stripe[3233] = 24'hffffff;
assign target_only_stripe[3234] = 24'hffffff;
assign target_only_stripe[3235] = 24'hffffff;
assign target_only_stripe[3236] = 24'hffffff;
assign target_only_stripe[3237] = 24'hffffff;
assign target_only_stripe[3238] = 24'hffffff;
assign target_only_stripe[3239] = 24'hffffff;
assign target_only_stripe[3240] = 24'hffffff;
assign target_only_stripe[3241] = 24'hffffff;
assign target_only_stripe[3242] = 24'hffffff;
assign target_only_stripe[3243] = 24'hffffff;
assign target_only_stripe[3244] = 24'hffffff;
assign target_only_stripe[3245] = 24'hffffff;
assign target_only_stripe[3246] = 24'hffffff;
assign target_only_stripe[3247] = 24'hffffff;
assign target_only_stripe[3248] = 24'hffffff;
assign target_only_stripe[3249] = 24'hffffff;
assign target_only_stripe[3250] = 24'hffffff;
assign target_only_stripe[3251] = 24'hffffff;
assign target_only_stripe[3252] = 24'hffffff;
assign target_only_stripe[3253] = 24'hffffff;
assign target_only_stripe[3254] = 24'hffffff;
assign target_only_stripe[3255] = 24'hffffff;
assign target_only_stripe[3256] = 24'hffffff;
assign target_only_stripe[3257] = 24'hd1b9ac;
assign target_only_stripe[3258] = 24'h1b1b1b;
assign target_only_stripe[3259] = 24'h000000;
assign target_only_stripe[3260] = 24'h000000;
assign target_only_stripe[3261] = 24'h000000;
assign target_only_stripe[3262] = 24'h000000;
assign target_only_stripe[3263] = 24'h000000;
assign target_only_stripe[3264] = 24'h000000;
assign target_only_stripe[3265] = 24'h000000;
assign target_only_stripe[3266] = 24'h000000;
assign target_only_stripe[3267] = 24'h000000;
assign target_only_stripe[3268] = 24'h000000;
assign target_only_stripe[3269] = 24'h000000;
assign target_only_stripe[3270] = 24'h000000;
assign target_only_stripe[3271] = 24'h000000;
assign target_only_stripe[3272] = 24'h000000;
assign target_only_stripe[3273] = 24'h000000;
assign target_only_stripe[3274] = 24'h000000;
assign target_only_stripe[3275] = 24'h000000;
assign target_only_stripe[3276] = 24'h000000;
assign target_only_stripe[3277] = 24'h000000;
assign target_only_stripe[3278] = 24'h000000;
assign target_only_stripe[3279] = 24'h000000;
assign target_only_stripe[3280] = 24'h000000;
assign target_only_stripe[3281] = 24'h000000;
assign target_only_stripe[3282] = 24'h000000;
assign target_only_stripe[3283] = 24'h000000;
assign target_only_stripe[3284] = 24'h000000;
assign target_only_stripe[3285] = 24'h000000;
assign target_only_stripe[3286] = 24'h000000;
assign target_only_stripe[3287] = 24'h000000;
assign target_only_stripe[3288] = 24'h000000;
assign target_only_stripe[3289] = 24'h000000;
assign target_only_stripe[3290] = 24'h000000;
assign target_only_stripe[3291] = 24'h000000;
assign target_only_stripe[3292] = 24'h000000;
assign target_only_stripe[3293] = 24'h000000;
assign target_only_stripe[3294] = 24'h000000;
assign target_only_stripe[3295] = 24'h000000;
assign target_only_stripe[3296] = 24'h000000;
assign target_only_stripe[3297] = 24'h000000;
assign target_only_stripe[3298] = 24'h000000;
assign target_only_stripe[3299] = 24'h000000;
assign target_only_stripe[3300] = 24'h000000;
assign target_only_stripe[3301] = 24'h000000;
assign target_only_stripe[3302] = 24'h000000;
assign target_only_stripe[3303] = 24'h000000;
assign target_only_stripe[3304] = 24'h000000;
assign target_only_stripe[3305] = 24'h000000;
assign target_only_stripe[3306] = 24'h000000;
assign target_only_stripe[3307] = 24'h000000;
assign target_only_stripe[3308] = 24'h000000;
assign target_only_stripe[3309] = 24'h000000;
assign target_only_stripe[3310] = 24'h000000;
assign target_only_stripe[3311] = 24'h000000;
assign target_only_stripe[3312] = 24'h000000;
assign target_only_stripe[3313] = 24'h000000;
assign target_only_stripe[3314] = 24'h000000;
assign target_only_stripe[3315] = 24'h000000;
assign target_only_stripe[3316] = 24'h000000;
assign target_only_stripe[3317] = 24'h000000;
assign target_only_stripe[3318] = 24'h000000;
assign target_only_stripe[3319] = 24'h000000;
assign target_only_stripe[3320] = 24'h000000;
assign target_only_stripe[3321] = 24'h121212;
assign target_only_stripe[3322] = 24'he8e6e6;
assign target_only_stripe[3323] = 24'hffffff;
assign target_only_stripe[3324] = 24'hffffff;
assign target_only_stripe[3325] = 24'hffffff;
assign target_only_stripe[3326] = 24'hffffff;
assign target_only_stripe[3327] = 24'hffffff;
assign target_only_stripe[3328] = 24'hffffff;
assign target_only_stripe[3329] = 24'hffffff;
assign target_only_stripe[3330] = 24'hffffff;
assign target_only_stripe[3331] = 24'hffffff;
assign target_only_stripe[3332] = 24'hffffff;
assign target_only_stripe[3333] = 24'hffffff;
assign target_only_stripe[3334] = 24'hffffff;
assign target_only_stripe[3335] = 24'hffffff;
assign target_only_stripe[3336] = 24'hffffff;
assign target_only_stripe[3337] = 24'hffffff;
assign target_only_stripe[3338] = 24'hffffff;
assign target_only_stripe[3339] = 24'hffffff;
assign target_only_stripe[3340] = 24'hffffff;
assign target_only_stripe[3341] = 24'hffffff;
assign target_only_stripe[3342] = 24'hffffff;
assign target_only_stripe[3343] = 24'hffffff;
assign target_only_stripe[3344] = 24'hffffff;
assign target_only_stripe[3345] = 24'hffffff;
assign target_only_stripe[3346] = 24'hffffff;
assign target_only_stripe[3347] = 24'hffffff;
assign target_only_stripe[3348] = 24'hffffff;
assign target_only_stripe[3349] = 24'hffffff;
assign target_only_stripe[3350] = 24'hffffff;
assign target_only_stripe[3351] = 24'hf4eae1;
assign target_only_stripe[3352] = 24'hffffff;
assign target_only_stripe[3353] = 24'hf0e8de;
assign target_only_stripe[3354] = 24'hffffff;
assign target_only_stripe[3355] = 24'hbebebe;
assign target_only_stripe[3356] = 24'h000000;
assign target_only_stripe[3357] = 24'h000000;
assign target_only_stripe[3358] = 24'h000000;
assign target_only_stripe[3359] = 24'h000000;
assign target_only_stripe[3360] = 24'h000000;
assign target_only_stripe[3361] = 24'h000000;
assign target_only_stripe[3362] = 24'h000000;
assign target_only_stripe[3363] = 24'h000000;
assign target_only_stripe[3364] = 24'h000000;
assign target_only_stripe[3365] = 24'h000000;
assign target_only_stripe[3366] = 24'h000000;
assign target_only_stripe[3367] = 24'h000000;
assign target_only_stripe[3368] = 24'h000000;
assign target_only_stripe[3369] = 24'h000000;
assign target_only_stripe[3370] = 24'h000000;
assign target_only_stripe[3371] = 24'h000000;
assign target_only_stripe[3372] = 24'h000000;
assign target_only_stripe[3373] = 24'h000000;
assign target_only_stripe[3374] = 24'h000000;
assign target_only_stripe[3375] = 24'h000000;
assign target_only_stripe[3376] = 24'h000000;
assign target_only_stripe[3377] = 24'h000000;
assign target_only_stripe[3378] = 24'h000000;
assign target_only_stripe[3379] = 24'h000000;
assign target_only_stripe[3380] = 24'h000000;
assign target_only_stripe[3381] = 24'h000000;
assign target_only_stripe[3382] = 24'h000000;
assign target_only_stripe[3383] = 24'h000000;
assign target_only_stripe[3384] = 24'h000000;
assign target_only_stripe[3385] = 24'h000000;
assign target_only_stripe[3386] = 24'h000000;
assign target_only_stripe[3387] = 24'h000000;
assign target_only_stripe[3388] = 24'ha3a3a3;
assign target_only_stripe[3389] = 24'hffffff;
assign target_only_stripe[3390] = 24'hffffff;
assign target_only_stripe[3391] = 24'hffffff;
assign target_only_stripe[3392] = 24'hffffff;
assign target_only_stripe[3393] = 24'hffffff;
assign target_only_stripe[3394] = 24'hffffff;
assign target_only_stripe[3395] = 24'hffffff;
assign target_only_stripe[3396] = 24'hffffff;
assign target_only_stripe[3397] = 24'hffffff;
assign target_only_stripe[3398] = 24'hffffff;
assign target_only_stripe[3399] = 24'hffffff;
assign target_only_stripe[3400] = 24'hffffff;
assign target_only_stripe[3401] = 24'hffffff;
assign target_only_stripe[3402] = 24'hffffff;
assign target_only_stripe[3403] = 24'hffffff;
assign target_only_stripe[3404] = 24'hffffff;
assign target_only_stripe[3405] = 24'hffffff;
assign target_only_stripe[3406] = 24'hffffff;
assign target_only_stripe[3407] = 24'hffffff;
assign target_only_stripe[3408] = 24'hffffff;
assign target_only_stripe[3409] = 24'hffffff;
assign target_only_stripe[3410] = 24'hffffff;
assign target_only_stripe[3411] = 24'hffffff;
assign target_only_stripe[3412] = 24'hffffff;
assign target_only_stripe[3413] = 24'hffffff;
assign target_only_stripe[3414] = 24'hffffff;
assign target_only_stripe[3415] = 24'hffffff;
assign target_only_stripe[3416] = 24'hffffff;
assign target_only_stripe[3417] = 24'hffffff;
assign target_only_stripe[3418] = 24'hffffff;
assign target_only_stripe[3419] = 24'hffffff;
assign target_only_stripe[3420] = 24'hffffff;
assign target_only_stripe[3421] = 24'hffffff;
assign target_only_stripe[3422] = 24'h383838;
assign target_only_stripe[3423] = 24'h000000;
assign target_only_stripe[3424] = 24'h000000;
assign target_only_stripe[3425] = 24'h000000;
assign target_only_stripe[3426] = 24'h000000;
assign target_only_stripe[3427] = 24'h000000;
assign target_only_stripe[3428] = 24'h000000;
assign target_only_stripe[3429] = 24'h000000;
assign target_only_stripe[3430] = 24'h000000;
assign target_only_stripe[3431] = 24'h000000;
assign target_only_stripe[3432] = 24'h000000;
assign target_only_stripe[3433] = 24'h000000;
assign target_only_stripe[3434] = 24'h000000;
assign target_only_stripe[3435] = 24'h000000;
assign target_only_stripe[3436] = 24'h000000;
assign target_only_stripe[3437] = 24'h000000;
assign target_only_stripe[3438] = 24'h000000;
assign target_only_stripe[3439] = 24'h000000;
assign target_only_stripe[3440] = 24'h000000;
assign target_only_stripe[3441] = 24'h000000;
assign target_only_stripe[3442] = 24'h000000;
assign target_only_stripe[3443] = 24'h000000;
assign target_only_stripe[3444] = 24'h000000;
assign target_only_stripe[3445] = 24'h000000;
assign target_only_stripe[3446] = 24'h000000;
assign target_only_stripe[3447] = 24'h000000;
assign target_only_stripe[3448] = 24'h000000;
assign target_only_stripe[3449] = 24'h000000;
assign target_only_stripe[3450] = 24'h000000;
assign target_only_stripe[3451] = 24'h000000;
assign target_only_stripe[3452] = 24'h000000;
assign target_only_stripe[3453] = 24'h000000;
assign target_only_stripe[3454] = 24'h000000;
assign target_only_stripe[3455] = 24'h000000;
assign target_only_stripe[3456] = 24'h000000;
assign target_only_stripe[3457] = 24'h000000;
assign target_only_stripe[3458] = 24'h000000;
assign target_only_stripe[3459] = 24'h000000;
assign target_only_stripe[3460] = 24'h000000;
assign target_only_stripe[3461] = 24'h000000;
assign target_only_stripe[3462] = 24'h000000;
assign target_only_stripe[3463] = 24'h000000;
assign target_only_stripe[3464] = 24'h000000;
assign target_only_stripe[3465] = 24'h000000;
assign target_only_stripe[3466] = 24'h000000;
assign target_only_stripe[3467] = 24'h000000;
assign target_only_stripe[3468] = 24'h000000;
assign target_only_stripe[3469] = 24'h000000;
assign target_only_stripe[3470] = 24'h000000;
assign target_only_stripe[3471] = 24'h000000;
assign target_only_stripe[3472] = 24'h000000;
assign target_only_stripe[3473] = 24'h000000;
assign target_only_stripe[3474] = 24'h000000;
assign target_only_stripe[3475] = 24'h000000;
assign target_only_stripe[3476] = 24'h000000;
assign target_only_stripe[3477] = 24'h000000;
assign target_only_stripe[3478] = 24'h000000;
assign target_only_stripe[3479] = 24'h000000;
assign target_only_stripe[3480] = 24'h000000;
assign target_only_stripe[3481] = 24'h000000;
assign target_only_stripe[3482] = 24'h000000;
assign target_only_stripe[3483] = 24'h000000;
assign target_only_stripe[3484] = 24'h000000;
assign target_only_stripe[3485] = 24'h000000;
assign target_only_stripe[3486] = 24'h313131;
assign target_only_stripe[3487] = 24'hffffff;
assign target_only_stripe[3488] = 24'hffffff;
assign target_only_stripe[3489] = 24'hffffff;
assign target_only_stripe[3490] = 24'hffffff;
assign target_only_stripe[3491] = 24'hffffff;
assign target_only_stripe[3492] = 24'hffffff;
assign target_only_stripe[3493] = 24'hffffff;
assign target_only_stripe[3494] = 24'hffffff;
assign target_only_stripe[3495] = 24'hffffff;
assign target_only_stripe[3496] = 24'hffffff;
assign target_only_stripe[3497] = 24'hffffff;
assign target_only_stripe[3498] = 24'hffffff;
assign target_only_stripe[3499] = 24'hffffff;
assign target_only_stripe[3500] = 24'hffffff;
assign target_only_stripe[3501] = 24'hffffff;
assign target_only_stripe[3502] = 24'hffffff;
assign target_only_stripe[3503] = 24'hffffff;
assign target_only_stripe[3504] = 24'hffffff;
assign target_only_stripe[3505] = 24'hffffff;
assign target_only_stripe[3506] = 24'hffffff;
assign target_only_stripe[3507] = 24'hffffff;
assign target_only_stripe[3508] = 24'hffffff;
assign target_only_stripe[3509] = 24'hffffff;
assign target_only_stripe[3510] = 24'hffffff;
assign target_only_stripe[3511] = 24'hffffff;
assign target_only_stripe[3512] = 24'hffffff;
assign target_only_stripe[3513] = 24'hffffff;
assign target_only_stripe[3514] = 24'hffffff;
assign target_only_stripe[3515] = 24'hffffff;
assign target_only_stripe[3516] = 24'hffffff;
assign target_only_stripe[3517] = 24'hffffff;
assign target_only_stripe[3518] = 24'hffffff;
assign target_only_stripe[3519] = 24'hffffff;
assign target_only_stripe[3520] = 24'haaaaaa;
assign target_only_stripe[3521] = 24'h000000;
assign target_only_stripe[3522] = 24'h000000;
assign target_only_stripe[3523] = 24'h000000;
assign target_only_stripe[3524] = 24'h000000;
assign target_only_stripe[3525] = 24'h000000;
assign target_only_stripe[3526] = 24'h000000;
assign target_only_stripe[3527] = 24'h000000;
assign target_only_stripe[3528] = 24'h000000;
assign target_only_stripe[3529] = 24'h000000;
assign target_only_stripe[3530] = 24'h000000;
assign target_only_stripe[3531] = 24'h000000;
assign target_only_stripe[3532] = 24'h000000;
assign target_only_stripe[3533] = 24'h000000;
assign target_only_stripe[3534] = 24'h000000;
assign target_only_stripe[3535] = 24'h000000;
assign target_only_stripe[3536] = 24'h000000;
assign target_only_stripe[3537] = 24'h000000;
assign target_only_stripe[3538] = 24'h000000;
assign target_only_stripe[3539] = 24'h000000;
assign target_only_stripe[3540] = 24'h000000;
assign target_only_stripe[3541] = 24'h000000;
assign target_only_stripe[3542] = 24'h000000;
assign target_only_stripe[3543] = 24'h000000;
assign target_only_stripe[3544] = 24'h000000;
assign target_only_stripe[3545] = 24'h000000;
assign target_only_stripe[3546] = 24'h000000;
assign target_only_stripe[3547] = 24'h000000;
assign target_only_stripe[3548] = 24'h000000;
assign target_only_stripe[3549] = 24'h000000;
assign target_only_stripe[3550] = 24'h000000;
assign target_only_stripe[3551] = 24'h000000;
assign target_only_stripe[3552] = 24'h000000;
assign target_only_stripe[3553] = 24'hd7d7d7;
assign target_only_stripe[3554] = 24'hffffff;
assign target_only_stripe[3555] = 24'hffffff;
assign target_only_stripe[3556] = 24'hffffff;
assign target_only_stripe[3557] = 24'hffffff;
assign target_only_stripe[3558] = 24'hffffff;
assign target_only_stripe[3559] = 24'hffffff;
assign target_only_stripe[3560] = 24'hffffff;
assign target_only_stripe[3561] = 24'hffffff;
assign target_only_stripe[3562] = 24'hffffff;
assign target_only_stripe[3563] = 24'hffffff;
assign target_only_stripe[3564] = 24'hffffff;
assign target_only_stripe[3565] = 24'hffffff;
assign target_only_stripe[3566] = 24'hffffff;
assign target_only_stripe[3567] = 24'hffffff;
assign target_only_stripe[3568] = 24'hffffff;
assign target_only_stripe[3569] = 24'hffffff;
assign target_only_stripe[3570] = 24'hffffff;
assign target_only_stripe[3571] = 24'hffffff;
assign target_only_stripe[3572] = 24'hffffff;
assign target_only_stripe[3573] = 24'hffffff;
assign target_only_stripe[3574] = 24'hffffff;
assign target_only_stripe[3575] = 24'hffffff;
assign target_only_stripe[3576] = 24'hffffff;
assign target_only_stripe[3577] = 24'hffffff;
assign target_only_stripe[3578] = 24'hffffff;
assign target_only_stripe[3579] = 24'hffffff;
assign target_only_stripe[3580] = 24'hffffff;
assign target_only_stripe[3581] = 24'hffffff;
assign target_only_stripe[3582] = 24'hffffff;
assign target_only_stripe[3583] = 24'hffffff;
assign target_only_stripe[3584] = 24'hffffff;
assign target_only_stripe[3585] = 24'hffffff;
assign target_only_stripe[3586] = 24'hddc0b0;
assign target_only_stripe[3587] = 24'h1b1b1b;
assign target_only_stripe[3588] = 24'h000000;
assign target_only_stripe[3589] = 24'h000000;
assign target_only_stripe[3590] = 24'h000000;
assign target_only_stripe[3591] = 24'h000000;
assign target_only_stripe[3592] = 24'h000000;
assign target_only_stripe[3593] = 24'h000000;
assign target_only_stripe[3594] = 24'h000000;
assign target_only_stripe[3595] = 24'h000000;
assign target_only_stripe[3596] = 24'h000000;
assign target_only_stripe[3597] = 24'h000000;
assign target_only_stripe[3598] = 24'h000000;
assign target_only_stripe[3599] = 24'h000000;
assign target_only_stripe[3600] = 24'h000000;
assign target_only_stripe[3601] = 24'h000000;
assign target_only_stripe[3602] = 24'h000000;
assign target_only_stripe[3603] = 24'h000000;
assign target_only_stripe[3604] = 24'h000000;
assign target_only_stripe[3605] = 24'h000000;
assign target_only_stripe[3606] = 24'h000000;
assign target_only_stripe[3607] = 24'h000000;
assign target_only_stripe[3608] = 24'h000000;
assign target_only_stripe[3609] = 24'h000000;
assign target_only_stripe[3610] = 24'h000000;
assign target_only_stripe[3611] = 24'h000000;
assign target_only_stripe[3612] = 24'h000000;
assign target_only_stripe[3613] = 24'h000000;
assign target_only_stripe[3614] = 24'h000000;
assign target_only_stripe[3615] = 24'h000000;
assign target_only_stripe[3616] = 24'h000000;
assign target_only_stripe[3617] = 24'h000000;
assign target_only_stripe[3618] = 24'h000000;
assign target_only_stripe[3619] = 24'h000000;
assign target_only_stripe[3620] = 24'h000000;
assign target_only_stripe[3621] = 24'h000000;
assign target_only_stripe[3622] = 24'h000000;
assign target_only_stripe[3623] = 24'h000000;
assign target_only_stripe[3624] = 24'h000000;
assign target_only_stripe[3625] = 24'h000000;
assign target_only_stripe[3626] = 24'h000000;
assign target_only_stripe[3627] = 24'h000000;
assign target_only_stripe[3628] = 24'h000000;
assign target_only_stripe[3629] = 24'h000000;
assign target_only_stripe[3630] = 24'h000000;
assign target_only_stripe[3631] = 24'h000000;
assign target_only_stripe[3632] = 24'h000000;
assign target_only_stripe[3633] = 24'h000000;
assign target_only_stripe[3634] = 24'h000000;
assign target_only_stripe[3635] = 24'h000000;
assign target_only_stripe[3636] = 24'h000000;
assign target_only_stripe[3637] = 24'h000000;
assign target_only_stripe[3638] = 24'h000000;
assign target_only_stripe[3639] = 24'h000000;
assign target_only_stripe[3640] = 24'h000000;
assign target_only_stripe[3641] = 24'h000000;
assign target_only_stripe[3642] = 24'h000000;
assign target_only_stripe[3643] = 24'h000000;
assign target_only_stripe[3644] = 24'h000000;
assign target_only_stripe[3645] = 24'h000000;
assign target_only_stripe[3646] = 24'h000000;
assign target_only_stripe[3647] = 24'h000000;
assign target_only_stripe[3648] = 24'h000000;
assign target_only_stripe[3649] = 24'h000000;
assign target_only_stripe[3650] = 24'h121212;
assign target_only_stripe[3651] = 24'he8e6e6;
assign target_only_stripe[3652] = 24'hffffff;
assign target_only_stripe[3653] = 24'hffffff;
assign target_only_stripe[3654] = 24'hffffff;
assign target_only_stripe[3655] = 24'hffffff;
assign target_only_stripe[3656] = 24'hffffff;
assign target_only_stripe[3657] = 24'hffffff;
assign target_only_stripe[3658] = 24'hffffff;
assign target_only_stripe[3659] = 24'hffffff;
assign target_only_stripe[3660] = 24'hffffff;
assign target_only_stripe[3661] = 24'hffffff;
assign target_only_stripe[3662] = 24'hffffff;
assign target_only_stripe[3663] = 24'hffffff;
assign target_only_stripe[3664] = 24'hffffff;
assign target_only_stripe[3665] = 24'hffffff;
assign target_only_stripe[3666] = 24'hffffff;
assign target_only_stripe[3667] = 24'hffffff;
assign target_only_stripe[3668] = 24'hffffff;
assign target_only_stripe[3669] = 24'hffffff;
assign target_only_stripe[3670] = 24'hffffff;
assign target_only_stripe[3671] = 24'hffffff;
assign target_only_stripe[3672] = 24'hffffff;
assign target_only_stripe[3673] = 24'hffffff;
assign target_only_stripe[3674] = 24'hffffff;
assign target_only_stripe[3675] = 24'hffffff;
assign target_only_stripe[3676] = 24'hffffff;
assign target_only_stripe[3677] = 24'hffffff;
assign target_only_stripe[3678] = 24'hffffff;
assign target_only_stripe[3679] = 24'hffffff;
assign target_only_stripe[3680] = 24'hf9f5f2;
assign target_only_stripe[3681] = 24'hffffff;
assign target_only_stripe[3682] = 24'hfaf7f5;
assign target_only_stripe[3683] = 24'hffffff;
assign target_only_stripe[3684] = 24'hc9c9c9;
assign target_only_stripe[3685] = 24'h000000;
assign target_only_stripe[3686] = 24'h000000;
assign target_only_stripe[3687] = 24'h000000;
assign target_only_stripe[3688] = 24'h000000;
assign target_only_stripe[3689] = 24'h000000;
assign target_only_stripe[3690] = 24'h000000;
assign target_only_stripe[3691] = 24'h000000;
assign target_only_stripe[3692] = 24'h000000;
assign target_only_stripe[3693] = 24'h000000;
assign target_only_stripe[3694] = 24'h000000;
assign target_only_stripe[3695] = 24'h000000;
assign target_only_stripe[3696] = 24'h000000;
assign target_only_stripe[3697] = 24'h000000;
assign target_only_stripe[3698] = 24'h000000;
assign target_only_stripe[3699] = 24'h000000;
assign target_only_stripe[3700] = 24'h000000;
assign target_only_stripe[3701] = 24'h000000;
assign target_only_stripe[3702] = 24'h000000;
assign target_only_stripe[3703] = 24'h000000;
assign target_only_stripe[3704] = 24'h000000;
assign target_only_stripe[3705] = 24'h000000;
assign target_only_stripe[3706] = 24'h000000;
assign target_only_stripe[3707] = 24'h000000;
assign target_only_stripe[3708] = 24'h000000;
assign target_only_stripe[3709] = 24'h000000;
assign target_only_stripe[3710] = 24'h000000;
assign target_only_stripe[3711] = 24'h000000;
assign target_only_stripe[3712] = 24'h000000;
assign target_only_stripe[3713] = 24'h000000;
assign target_only_stripe[3714] = 24'h000000;
assign target_only_stripe[3715] = 24'h000000;
assign target_only_stripe[3716] = 24'h000000;
assign target_only_stripe[3717] = 24'hb8b8b8;
assign target_only_stripe[3718] = 24'hffffff;
assign target_only_stripe[3719] = 24'hffffff;
assign target_only_stripe[3720] = 24'hffffff;
assign target_only_stripe[3721] = 24'hffffff;
assign target_only_stripe[3722] = 24'hffffff;
assign target_only_stripe[3723] = 24'hffffff;
assign target_only_stripe[3724] = 24'hffffff;
assign target_only_stripe[3725] = 24'hffffff;
assign target_only_stripe[3726] = 24'hffffff;
assign target_only_stripe[3727] = 24'hffffff;
assign target_only_stripe[3728] = 24'hffffff;
assign target_only_stripe[3729] = 24'hffffff;
assign target_only_stripe[3730] = 24'hffffff;
assign target_only_stripe[3731] = 24'hffffff;
assign target_only_stripe[3732] = 24'hffffff;
assign target_only_stripe[3733] = 24'hffffff;
assign target_only_stripe[3734] = 24'hffffff;
assign target_only_stripe[3735] = 24'hffffff;
assign target_only_stripe[3736] = 24'hffffff;
assign target_only_stripe[3737] = 24'hffffff;
assign target_only_stripe[3738] = 24'hffffff;
assign target_only_stripe[3739] = 24'hffffff;
assign target_only_stripe[3740] = 24'hffffff;
assign target_only_stripe[3741] = 24'hffffff;
assign target_only_stripe[3742] = 24'hffffff;
assign target_only_stripe[3743] = 24'hffffff;
assign target_only_stripe[3744] = 24'hffffff;
assign target_only_stripe[3745] = 24'hffffff;
assign target_only_stripe[3746] = 24'hffffff;
assign target_only_stripe[3747] = 24'hffffff;
assign target_only_stripe[3748] = 24'hffffff;
assign target_only_stripe[3749] = 24'hffffff;
assign target_only_stripe[3750] = 24'hffffff;
assign target_only_stripe[3751] = 24'h282828;
assign target_only_stripe[3752] = 24'h000000;
assign target_only_stripe[3753] = 24'h000000;
assign target_only_stripe[3754] = 24'h000000;
assign target_only_stripe[3755] = 24'h000000;
assign target_only_stripe[3756] = 24'h000000;
assign target_only_stripe[3757] = 24'h000000;
assign target_only_stripe[3758] = 24'h000000;
assign target_only_stripe[3759] = 24'h000000;
assign target_only_stripe[3760] = 24'h000000;
assign target_only_stripe[3761] = 24'h000000;
assign target_only_stripe[3762] = 24'h000000;
assign target_only_stripe[3763] = 24'h000000;
assign target_only_stripe[3764] = 24'h000000;
assign target_only_stripe[3765] = 24'h000000;
assign target_only_stripe[3766] = 24'h000000;
assign target_only_stripe[3767] = 24'h000000;
assign target_only_stripe[3768] = 24'h000000;
assign target_only_stripe[3769] = 24'h000000;
assign target_only_stripe[3770] = 24'h000000;
assign target_only_stripe[3771] = 24'h000000;
assign target_only_stripe[3772] = 24'h000000;
assign target_only_stripe[3773] = 24'h000000;
assign target_only_stripe[3774] = 24'h000000;
assign target_only_stripe[3775] = 24'h000000;
assign target_only_stripe[3776] = 24'h000000;
assign target_only_stripe[3777] = 24'h000000;
assign target_only_stripe[3778] = 24'h000000;
assign target_only_stripe[3779] = 24'h000000;
assign target_only_stripe[3780] = 24'h000000;
assign target_only_stripe[3781] = 24'h000000;
assign target_only_stripe[3782] = 24'h000000;
assign target_only_stripe[3783] = 24'h000000;
assign target_only_stripe[3784] = 24'h000000;
assign target_only_stripe[3785] = 24'h000000;
assign target_only_stripe[3786] = 24'h000000;
assign target_only_stripe[3787] = 24'h000000;
assign target_only_stripe[3788] = 24'h000000;
assign target_only_stripe[3789] = 24'h000000;
assign target_only_stripe[3790] = 24'h000000;
assign target_only_stripe[3791] = 24'h000000;
assign target_only_stripe[3792] = 24'h000000;
assign target_only_stripe[3793] = 24'h000000;
assign target_only_stripe[3794] = 24'h000000;
assign target_only_stripe[3795] = 24'h000000;
assign target_only_stripe[3796] = 24'h000000;
assign target_only_stripe[3797] = 24'h000000;
assign target_only_stripe[3798] = 24'h000000;
assign target_only_stripe[3799] = 24'h000000;
assign target_only_stripe[3800] = 24'h000000;
assign target_only_stripe[3801] = 24'h000000;
assign target_only_stripe[3802] = 24'h000000;
assign target_only_stripe[3803] = 24'h000000;
assign target_only_stripe[3804] = 24'h000000;
assign target_only_stripe[3805] = 24'h000000;
assign target_only_stripe[3806] = 24'h000000;
assign target_only_stripe[3807] = 24'h000000;
assign target_only_stripe[3808] = 24'h000000;
assign target_only_stripe[3809] = 24'h000000;
assign target_only_stripe[3810] = 24'h000000;
assign target_only_stripe[3811] = 24'h000000;
assign target_only_stripe[3812] = 24'h000000;
assign target_only_stripe[3813] = 24'h000000;
assign target_only_stripe[3814] = 24'h000000;
assign target_only_stripe[3815] = 24'h222222;
assign target_only_stripe[3816] = 24'hffffff;
assign target_only_stripe[3817] = 24'hffffff;
assign target_only_stripe[3818] = 24'hffffff;
assign target_only_stripe[3819] = 24'hffffff;
assign target_only_stripe[3820] = 24'hffffff;
assign target_only_stripe[3821] = 24'hffffff;
assign target_only_stripe[3822] = 24'hffffff;
assign target_only_stripe[3823] = 24'hffffff;
assign target_only_stripe[3824] = 24'hffffff;
assign target_only_stripe[3825] = 24'hffffff;
assign target_only_stripe[3826] = 24'hffffff;
assign target_only_stripe[3827] = 24'hffffff;
assign target_only_stripe[3828] = 24'hffffff;
assign target_only_stripe[3829] = 24'hffffff;
assign target_only_stripe[3830] = 24'hffffff;
assign target_only_stripe[3831] = 24'hffffff;
assign target_only_stripe[3832] = 24'hffffff;
assign target_only_stripe[3833] = 24'hffffff;
assign target_only_stripe[3834] = 24'hffffff;
assign target_only_stripe[3835] = 24'hffffff;
assign target_only_stripe[3836] = 24'hffffff;
assign target_only_stripe[3837] = 24'hffffff;
assign target_only_stripe[3838] = 24'hffffff;
assign target_only_stripe[3839] = 24'hffffff;
assign target_only_stripe[3840] = 24'hffffff;
assign target_only_stripe[3841] = 24'hffffff;
assign target_only_stripe[3842] = 24'hffffff;
assign target_only_stripe[3843] = 24'hffffff;
assign target_only_stripe[3844] = 24'hffffff;
assign target_only_stripe[3845] = 24'hffffff;
assign target_only_stripe[3846] = 24'hffffff;
assign target_only_stripe[3847] = 24'hffffff;
assign target_only_stripe[3848] = 24'hffffff;
assign target_only_stripe[3849] = 24'hd1d1d1;
assign target_only_stripe[3850] = 24'h000000;
assign target_only_stripe[3851] = 24'h000000;
assign target_only_stripe[3852] = 24'h000000;
assign target_only_stripe[3853] = 24'h000000;
assign target_only_stripe[3854] = 24'h000000;
assign target_only_stripe[3855] = 24'h000000;
assign target_only_stripe[3856] = 24'h000000;
assign target_only_stripe[3857] = 24'h000000;
assign target_only_stripe[3858] = 24'h000000;
assign target_only_stripe[3859] = 24'h000000;
assign target_only_stripe[3860] = 24'h000000;
assign target_only_stripe[3861] = 24'h000000;
assign target_only_stripe[3862] = 24'h000000;
assign target_only_stripe[3863] = 24'h000000;
assign target_only_stripe[3864] = 24'h000000;
assign target_only_stripe[3865] = 24'h000000;
assign target_only_stripe[3866] = 24'h000000;
assign target_only_stripe[3867] = 24'h000000;
assign target_only_stripe[3868] = 24'h000000;
assign target_only_stripe[3869] = 24'h000000;
assign target_only_stripe[3870] = 24'h000000;
assign target_only_stripe[3871] = 24'h000000;
assign target_only_stripe[3872] = 24'h000000;
assign target_only_stripe[3873] = 24'h000000;
assign target_only_stripe[3874] = 24'h000000;
assign target_only_stripe[3875] = 24'h000000;
assign target_only_stripe[3876] = 24'h000000;
assign target_only_stripe[3877] = 24'h000000;
assign target_only_stripe[3878] = 24'h000000;
assign target_only_stripe[3879] = 24'h000000;
assign target_only_stripe[3880] = 24'h000000;
assign target_only_stripe[3881] = 24'h000000;
assign target_only_stripe[3882] = 24'he1e1e1;
assign target_only_stripe[3883] = 24'hffffff;
assign target_only_stripe[3884] = 24'hffffff;
assign target_only_stripe[3885] = 24'hffffff;
assign target_only_stripe[3886] = 24'hffffff;
assign target_only_stripe[3887] = 24'hffffff;
assign target_only_stripe[3888] = 24'hffffff;
assign target_only_stripe[3889] = 24'hffffff;
assign target_only_stripe[3890] = 24'hffffff;
assign target_only_stripe[3891] = 24'hffffff;
assign target_only_stripe[3892] = 24'hffffff;
assign target_only_stripe[3893] = 24'hffffff;
assign target_only_stripe[3894] = 24'hffffff;
assign target_only_stripe[3895] = 24'hffffff;
assign target_only_stripe[3896] = 24'hffffff;
assign target_only_stripe[3897] = 24'hffffff;
assign target_only_stripe[3898] = 24'hffffff;
assign target_only_stripe[3899] = 24'hffffff;
assign target_only_stripe[3900] = 24'hffffff;
assign target_only_stripe[3901] = 24'hffffff;
assign target_only_stripe[3902] = 24'hffffff;
assign target_only_stripe[3903] = 24'hffffff;
assign target_only_stripe[3904] = 24'hffffff;
assign target_only_stripe[3905] = 24'hffffff;
assign target_only_stripe[3906] = 24'hffffff;
assign target_only_stripe[3907] = 24'hffffff;
assign target_only_stripe[3908] = 24'hffffff;
assign target_only_stripe[3909] = 24'hffffff;
assign target_only_stripe[3910] = 24'hffffff;
assign target_only_stripe[3911] = 24'hffffff;
assign target_only_stripe[3912] = 24'hffffff;
assign target_only_stripe[3913] = 24'hffffff;
assign target_only_stripe[3914] = 24'hffffff;
assign target_only_stripe[3915] = 24'hd9c0ae;
assign target_only_stripe[3916] = 24'h1b1b1b;
assign target_only_stripe[3917] = 24'h000000;
assign target_only_stripe[3918] = 24'h000000;
assign target_only_stripe[3919] = 24'h000000;
assign target_only_stripe[3920] = 24'h000000;
assign target_only_stripe[3921] = 24'h000000;
assign target_only_stripe[3922] = 24'h000000;
assign target_only_stripe[3923] = 24'h000000;
assign target_only_stripe[3924] = 24'h000000;
assign target_only_stripe[3925] = 24'h000000;
assign target_only_stripe[3926] = 24'h000000;
assign target_only_stripe[3927] = 24'h000000;
assign target_only_stripe[3928] = 24'h000000;
assign target_only_stripe[3929] = 24'h000000;
assign target_only_stripe[3930] = 24'h000000;
assign target_only_stripe[3931] = 24'h000000;
assign target_only_stripe[3932] = 24'h000000;
assign target_only_stripe[3933] = 24'h000000;
assign target_only_stripe[3934] = 24'h000000;
assign target_only_stripe[3935] = 24'h000000;
assign target_only_stripe[3936] = 24'h000000;
assign target_only_stripe[3937] = 24'h000000;
assign target_only_stripe[3938] = 24'h000000;
assign target_only_stripe[3939] = 24'h000000;
assign target_only_stripe[3940] = 24'h000000;
assign target_only_stripe[3941] = 24'h000000;
assign target_only_stripe[3942] = 24'h000000;
assign target_only_stripe[3943] = 24'h000000;
assign target_only_stripe[3944] = 24'h000000;
assign target_only_stripe[3945] = 24'h000000;
assign target_only_stripe[3946] = 24'h000000;
assign target_only_stripe[3947] = 24'h000000;
assign target_only_stripe[3948] = 24'h000000;
assign target_only_stripe[3949] = 24'h000000;
assign target_only_stripe[3950] = 24'h000000;
assign target_only_stripe[3951] = 24'h000000;
assign target_only_stripe[3952] = 24'h000000;
assign target_only_stripe[3953] = 24'h000000;
assign target_only_stripe[3954] = 24'h000000;
assign target_only_stripe[3955] = 24'h000000;
assign target_only_stripe[3956] = 24'h000000;
assign target_only_stripe[3957] = 24'h000000;
assign target_only_stripe[3958] = 24'h000000;
assign target_only_stripe[3959] = 24'h000000;
assign target_only_stripe[3960] = 24'h000000;
assign target_only_stripe[3961] = 24'h000000;
assign target_only_stripe[3962] = 24'h000000;
assign target_only_stripe[3963] = 24'h000000;
assign target_only_stripe[3964] = 24'h000000;
assign target_only_stripe[3965] = 24'h000000;
assign target_only_stripe[3966] = 24'h000000;
assign target_only_stripe[3967] = 24'h000000;
assign target_only_stripe[3968] = 24'h000000;
assign target_only_stripe[3969] = 24'h000000;
assign target_only_stripe[3970] = 24'h000000;
assign target_only_stripe[3971] = 24'h000000;
assign target_only_stripe[3972] = 24'h000000;
assign target_only_stripe[3973] = 24'h000000;
assign target_only_stripe[3974] = 24'h000000;
assign target_only_stripe[3975] = 24'h000000;
assign target_only_stripe[3976] = 24'h000000;
assign target_only_stripe[3977] = 24'h000000;
assign target_only_stripe[3978] = 24'h000000;
assign target_only_stripe[3979] = 24'h121212;
assign target_only_stripe[3980] = 24'he8e6e6;
assign target_only_stripe[3981] = 24'hffffff;
assign target_only_stripe[3982] = 24'hffffff;
assign target_only_stripe[3983] = 24'hffffff;
assign target_only_stripe[3984] = 24'hffffff;
assign target_only_stripe[3985] = 24'hffffff;
assign target_only_stripe[3986] = 24'hffffff;
assign target_only_stripe[3987] = 24'hffffff;
assign target_only_stripe[3988] = 24'hffffff;
assign target_only_stripe[3989] = 24'hffffff;
assign target_only_stripe[3990] = 24'hffffff;
assign target_only_stripe[3991] = 24'hffffff;
assign target_only_stripe[3992] = 24'hffffff;
assign target_only_stripe[3993] = 24'hffffff;
assign target_only_stripe[3994] = 24'hffffff;
assign target_only_stripe[3995] = 24'hffffff;
assign target_only_stripe[3996] = 24'hffffff;
assign target_only_stripe[3997] = 24'hffffff;
assign target_only_stripe[3998] = 24'hffffff;
assign target_only_stripe[3999] = 24'hffffff;
assign target_only_stripe[4000] = 24'hffffff;
assign target_only_stripe[4001] = 24'hffffff;
assign target_only_stripe[4002] = 24'hffffff;
assign target_only_stripe[4003] = 24'hffffff;
assign target_only_stripe[4004] = 24'hffffff;
assign target_only_stripe[4005] = 24'hffffff;
assign target_only_stripe[4006] = 24'hffffff;
assign target_only_stripe[4007] = 24'hffffff;
assign target_only_stripe[4008] = 24'hffffff;
assign target_only_stripe[4009] = 24'hffffff;
assign target_only_stripe[4010] = 24'hffffff;
assign target_only_stripe[4011] = 24'hffffff;
assign target_only_stripe[4012] = 24'hffffff;
assign target_only_stripe[4013] = 24'hc1c1c1;
assign target_only_stripe[4014] = 24'h000000;
assign target_only_stripe[4015] = 24'h000000;
assign target_only_stripe[4016] = 24'h000000;
assign target_only_stripe[4017] = 24'h000000;
assign target_only_stripe[4018] = 24'h000000;
assign target_only_stripe[4019] = 24'h000000;
assign target_only_stripe[4020] = 24'h000000;
assign target_only_stripe[4021] = 24'h000000;
assign target_only_stripe[4022] = 24'h000000;
assign target_only_stripe[4023] = 24'h000000;
assign target_only_stripe[4024] = 24'h000000;
assign target_only_stripe[4025] = 24'h000000;
assign target_only_stripe[4026] = 24'h000000;
assign target_only_stripe[4027] = 24'h000000;
assign target_only_stripe[4028] = 24'h000000;
assign target_only_stripe[4029] = 24'h000000;
assign target_only_stripe[4030] = 24'h000000;
assign target_only_stripe[4031] = 24'h000000;
assign target_only_stripe[4032] = 24'h000000;
assign target_only_stripe[4033] = 24'h000000;
assign target_only_stripe[4034] = 24'h000000;
assign target_only_stripe[4035] = 24'h000000;
assign target_only_stripe[4036] = 24'h000000;
assign target_only_stripe[4037] = 24'h000000;
assign target_only_stripe[4038] = 24'h000000;
assign target_only_stripe[4039] = 24'h000000;
assign target_only_stripe[4040] = 24'h000000;
assign target_only_stripe[4041] = 24'h000000;
assign target_only_stripe[4042] = 24'h000000;
assign target_only_stripe[4043] = 24'h000000;
assign target_only_stripe[4044] = 24'h000000;
assign target_only_stripe[4045] = 24'h000000;
assign target_only_stripe[4046] = 24'ha6a6a6;
assign target_only_stripe[4047] = 24'hffffff;
assign target_only_stripe[4048] = 24'hffffff;
assign target_only_stripe[4049] = 24'hffffff;
assign target_only_stripe[4050] = 24'hffffff;
assign target_only_stripe[4051] = 24'hffffff;
assign target_only_stripe[4052] = 24'hffffff;
assign target_only_stripe[4053] = 24'hffffff;
assign target_only_stripe[4054] = 24'hffffff;
assign target_only_stripe[4055] = 24'hffffff;
assign target_only_stripe[4056] = 24'hffffff;
assign target_only_stripe[4057] = 24'hffffff;
assign target_only_stripe[4058] = 24'hffffff;
assign target_only_stripe[4059] = 24'hffffff;
assign target_only_stripe[4060] = 24'hffffff;
assign target_only_stripe[4061] = 24'hffffff;
assign target_only_stripe[4062] = 24'hffffff;
assign target_only_stripe[4063] = 24'hffffff;
assign target_only_stripe[4064] = 24'hffffff;
assign target_only_stripe[4065] = 24'hffffff;
assign target_only_stripe[4066] = 24'hffffff;
assign target_only_stripe[4067] = 24'hffffff;
assign target_only_stripe[4068] = 24'hffffff;
assign target_only_stripe[4069] = 24'hffffff;
assign target_only_stripe[4070] = 24'hffffff;
assign target_only_stripe[4071] = 24'hffffff;
assign target_only_stripe[4072] = 24'hffffff;
assign target_only_stripe[4073] = 24'hffffff;
assign target_only_stripe[4074] = 24'hffffff;
assign target_only_stripe[4075] = 24'hffffff;
assign target_only_stripe[4076] = 24'hffffff;
assign target_only_stripe[4077] = 24'hffffff;
assign target_only_stripe[4078] = 24'hffffff;
assign target_only_stripe[4079] = 24'hffffff;
assign target_only_stripe[4080] = 24'h353535;
assign target_only_stripe[4081] = 24'h000000;
assign target_only_stripe[4082] = 24'h000000;
assign target_only_stripe[4083] = 24'h000000;
assign target_only_stripe[4084] = 24'h000000;
assign target_only_stripe[4085] = 24'h000000;
assign target_only_stripe[4086] = 24'h000000;
assign target_only_stripe[4087] = 24'h000000;
assign target_only_stripe[4088] = 24'h000000;
assign target_only_stripe[4089] = 24'h000000;
assign target_only_stripe[4090] = 24'h000000;
assign target_only_stripe[4091] = 24'h000000;
assign target_only_stripe[4092] = 24'h000000;
assign target_only_stripe[4093] = 24'h000000;
assign target_only_stripe[4094] = 24'h000000;
assign target_only_stripe[4095] = 24'h000000;
assign target_only_stripe[4096] = 24'h000000;
assign target_only_stripe[4097] = 24'h000000;
assign target_only_stripe[4098] = 24'h000000;
assign target_only_stripe[4099] = 24'h000000;
assign target_only_stripe[4100] = 24'h000000;
assign target_only_stripe[4101] = 24'h000000;
assign target_only_stripe[4102] = 24'h000000;
assign target_only_stripe[4103] = 24'h000000;
assign target_only_stripe[4104] = 24'h000000;
assign target_only_stripe[4105] = 24'h000000;
assign target_only_stripe[4106] = 24'h000000;
assign target_only_stripe[4107] = 24'h000000;
assign target_only_stripe[4108] = 24'h000000;
assign target_only_stripe[4109] = 24'h000000;
assign target_only_stripe[4110] = 24'h000000;
assign target_only_stripe[4111] = 24'h000000;
assign target_only_stripe[4112] = 24'h000000;
assign target_only_stripe[4113] = 24'h000000;
assign target_only_stripe[4114] = 24'h000000;
assign target_only_stripe[4115] = 24'h000000;
assign target_only_stripe[4116] = 24'h000000;
assign target_only_stripe[4117] = 24'h000000;
assign target_only_stripe[4118] = 24'h000000;
assign target_only_stripe[4119] = 24'h000000;
assign target_only_stripe[4120] = 24'h000000;
assign target_only_stripe[4121] = 24'h000000;
assign target_only_stripe[4122] = 24'h000000;
assign target_only_stripe[4123] = 24'h000000;
assign target_only_stripe[4124] = 24'h000000;
assign target_only_stripe[4125] = 24'h000000;
assign target_only_stripe[4126] = 24'h000000;
assign target_only_stripe[4127] = 24'h000000;
assign target_only_stripe[4128] = 24'h000000;
assign target_only_stripe[4129] = 24'h000000;
assign target_only_stripe[4130] = 24'h000000;
assign target_only_stripe[4131] = 24'h000000;
assign target_only_stripe[4132] = 24'h000000;
assign target_only_stripe[4133] = 24'h000000;
assign target_only_stripe[4134] = 24'h000000;
assign target_only_stripe[4135] = 24'h000000;
assign target_only_stripe[4136] = 24'h000000;
assign target_only_stripe[4137] = 24'h000000;
assign target_only_stripe[4138] = 24'h000000;
assign target_only_stripe[4139] = 24'h000000;
assign target_only_stripe[4140] = 24'h000000;
assign target_only_stripe[4141] = 24'h000000;
assign target_only_stripe[4142] = 24'h000000;
assign target_only_stripe[4143] = 24'h000000;
assign target_only_stripe[4144] = 24'h2e2e2e;
assign target_only_stripe[4145] = 24'hffffff;
assign target_only_stripe[4146] = 24'hffffff;
assign target_only_stripe[4147] = 24'hffffff;
assign target_only_stripe[4148] = 24'hffffff;
assign target_only_stripe[4149] = 24'hffffff;
assign target_only_stripe[4150] = 24'hffffff;
assign target_only_stripe[4151] = 24'hffffff;
assign target_only_stripe[4152] = 24'hffffff;
assign target_only_stripe[4153] = 24'hffffff;
assign target_only_stripe[4154] = 24'hffffff;
assign target_only_stripe[4155] = 24'hffffff;
assign target_only_stripe[4156] = 24'hffffff;
assign target_only_stripe[4157] = 24'hffffff;
assign target_only_stripe[4158] = 24'hffffff;
assign target_only_stripe[4159] = 24'hffffff;
assign target_only_stripe[4160] = 24'hffffff;
assign target_only_stripe[4161] = 24'hffffff;
assign target_only_stripe[4162] = 24'hffffff;
assign target_only_stripe[4163] = 24'hffffff;
assign target_only_stripe[4164] = 24'hffffff;
assign target_only_stripe[4165] = 24'hffffff;
assign target_only_stripe[4166] = 24'hffffff;
assign target_only_stripe[4167] = 24'hffffff;
assign target_only_stripe[4168] = 24'hffffff;
assign target_only_stripe[4169] = 24'hffffff;
assign target_only_stripe[4170] = 24'hffffff;
assign target_only_stripe[4171] = 24'hffffff;
assign target_only_stripe[4172] = 24'hffffff;
assign target_only_stripe[4173] = 24'hffffff;
assign target_only_stripe[4174] = 24'hffffff;
assign target_only_stripe[4175] = 24'hffffff;
assign target_only_stripe[4176] = 24'hffffff;
assign target_only_stripe[4177] = 24'hffffff;
assign target_only_stripe[4178] = 24'hadadad;
assign target_only_stripe[4179] = 24'h000000;
assign target_only_stripe[4180] = 24'h000000;
assign target_only_stripe[4181] = 24'h000000;
assign target_only_stripe[4182] = 24'h000000;
assign target_only_stripe[4183] = 24'h000000;
assign target_only_stripe[4184] = 24'h000000;
assign target_only_stripe[4185] = 24'h000000;
assign target_only_stripe[4186] = 24'h000000;
assign target_only_stripe[4187] = 24'h000000;
assign target_only_stripe[4188] = 24'h000000;
assign target_only_stripe[4189] = 24'h000000;
assign target_only_stripe[4190] = 24'h000000;
assign target_only_stripe[4191] = 24'h000000;
assign target_only_stripe[4192] = 24'h000000;
assign target_only_stripe[4193] = 24'h000000;
assign target_only_stripe[4194] = 24'h000000;
assign target_only_stripe[4195] = 24'h000000;
assign target_only_stripe[4196] = 24'h000000;
assign target_only_stripe[4197] = 24'h000000;
assign target_only_stripe[4198] = 24'h000000;
assign target_only_stripe[4199] = 24'h000000;
assign target_only_stripe[4200] = 24'h000000;
assign target_only_stripe[4201] = 24'h000000;
assign target_only_stripe[4202] = 24'h000000;
assign target_only_stripe[4203] = 24'h000000;
assign target_only_stripe[4204] = 24'h000000;
assign target_only_stripe[4205] = 24'h000000;
assign target_only_stripe[4206] = 24'h000000;
assign target_only_stripe[4207] = 24'h000000;
assign target_only_stripe[4208] = 24'h000000;
assign target_only_stripe[4209] = 24'h000000;
assign target_only_stripe[4210] = 24'h000000;
assign target_only_stripe[4211] = 24'hd9d9d9;
assign target_only_stripe[4212] = 24'hffffff;
assign target_only_stripe[4213] = 24'hffffff;
assign target_only_stripe[4214] = 24'hffffff;
assign target_only_stripe[4215] = 24'hffffff;
assign target_only_stripe[4216] = 24'hffffff;
assign target_only_stripe[4217] = 24'hffffff;
assign target_only_stripe[4218] = 24'hffffff;
assign target_only_stripe[4219] = 24'hffffff;
assign target_only_stripe[4220] = 24'hffffff;
assign target_only_stripe[4221] = 24'hffffff;
assign target_only_stripe[4222] = 24'hffffff;
assign target_only_stripe[4223] = 24'hffffff;
assign target_only_stripe[4224] = 24'hffffff;
assign target_only_stripe[4225] = 24'hffffff;
assign target_only_stripe[4226] = 24'hffffff;
assign target_only_stripe[4227] = 24'hffffff;
assign target_only_stripe[4228] = 24'hffffff;
assign target_only_stripe[4229] = 24'hffffff;
assign target_only_stripe[4230] = 24'hffffff;
assign target_only_stripe[4231] = 24'hffffff;
assign target_only_stripe[4232] = 24'hffffff;
assign target_only_stripe[4233] = 24'hffffff;
assign target_only_stripe[4234] = 24'hffffff;
assign target_only_stripe[4235] = 24'hffffff;
assign target_only_stripe[4236] = 24'hffffff;
assign target_only_stripe[4237] = 24'hffffff;
assign target_only_stripe[4238] = 24'hffffff;
assign target_only_stripe[4239] = 24'hffffff;
assign target_only_stripe[4240] = 24'hffffff;
assign target_only_stripe[4241] = 24'hffffff;
assign target_only_stripe[4242] = 24'hffffff;
assign target_only_stripe[4243] = 24'hffffff;
assign target_only_stripe[4244] = 24'hd5bdad;
assign target_only_stripe[4245] = 24'h1b1b1b;
assign target_only_stripe[4246] = 24'h000000;
assign target_only_stripe[4247] = 24'h000000;
assign target_only_stripe[4248] = 24'h000000;
assign target_only_stripe[4249] = 24'h000000;
assign target_only_stripe[4250] = 24'h000000;
assign target_only_stripe[4251] = 24'h000000;
assign target_only_stripe[4252] = 24'h000000;
assign target_only_stripe[4253] = 24'h000000;
assign target_only_stripe[4254] = 24'h000000;
assign target_only_stripe[4255] = 24'h000000;
assign target_only_stripe[4256] = 24'h000000;
assign target_only_stripe[4257] = 24'h000000;
assign target_only_stripe[4258] = 24'h000000;
assign target_only_stripe[4259] = 24'h000000;
assign target_only_stripe[4260] = 24'h000000;
assign target_only_stripe[4261] = 24'h000000;
assign target_only_stripe[4262] = 24'h000000;
assign target_only_stripe[4263] = 24'h000000;
assign target_only_stripe[4264] = 24'h000000;
assign target_only_stripe[4265] = 24'h000000;
assign target_only_stripe[4266] = 24'h000000;
assign target_only_stripe[4267] = 24'h000000;
assign target_only_stripe[4268] = 24'h000000;
assign target_only_stripe[4269] = 24'h000000;
assign target_only_stripe[4270] = 24'h000000;
assign target_only_stripe[4271] = 24'h000000;
assign target_only_stripe[4272] = 24'h000000;
assign target_only_stripe[4273] = 24'h000000;
assign target_only_stripe[4274] = 24'h000000;
assign target_only_stripe[4275] = 24'h000000;
assign target_only_stripe[4276] = 24'h000000;
assign target_only_stripe[4277] = 24'h000000;
assign target_only_stripe[4278] = 24'h000000;
assign target_only_stripe[4279] = 24'h000000;
assign target_only_stripe[4280] = 24'h000000;
assign target_only_stripe[4281] = 24'h000000;
assign target_only_stripe[4282] = 24'h000000;
assign target_only_stripe[4283] = 24'h000000;
assign target_only_stripe[4284] = 24'h000000;
assign target_only_stripe[4285] = 24'h000000;
assign target_only_stripe[4286] = 24'h000000;
assign target_only_stripe[4287] = 24'h000000;
assign target_only_stripe[4288] = 24'h000000;
assign target_only_stripe[4289] = 24'h000000;
assign target_only_stripe[4290] = 24'h000000;
assign target_only_stripe[4291] = 24'h000000;
assign target_only_stripe[4292] = 24'h000000;
assign target_only_stripe[4293] = 24'h000000;
assign target_only_stripe[4294] = 24'h000000;
assign target_only_stripe[4295] = 24'h000000;
assign target_only_stripe[4296] = 24'h000000;
assign target_only_stripe[4297] = 24'h000000;
assign target_only_stripe[4298] = 24'h000000;
assign target_only_stripe[4299] = 24'h000000;
assign target_only_stripe[4300] = 24'h000000;
assign target_only_stripe[4301] = 24'h000000;
assign target_only_stripe[4302] = 24'h000000;
assign target_only_stripe[4303] = 24'h000000;
assign target_only_stripe[4304] = 24'h000000;
assign target_only_stripe[4305] = 24'h000000;
assign target_only_stripe[4306] = 24'h000000;
assign target_only_stripe[4307] = 24'h000000;
assign target_only_stripe[4308] = 24'h121212;
assign target_only_stripe[4309] = 24'he8e6e6;
assign target_only_stripe[4310] = 24'hffffff;
assign target_only_stripe[4311] = 24'hffffff;
assign target_only_stripe[4312] = 24'hffffff;
assign target_only_stripe[4313] = 24'hffffff;
assign target_only_stripe[4314] = 24'hffffff;
assign target_only_stripe[4315] = 24'hffffff;
assign target_only_stripe[4316] = 24'hffffff;
assign target_only_stripe[4317] = 24'hffffff;
assign target_only_stripe[4318] = 24'hffffff;
assign target_only_stripe[4319] = 24'hffffff;
assign target_only_stripe[4320] = 24'hffffff;
assign target_only_stripe[4321] = 24'hffffff;
assign target_only_stripe[4322] = 24'hffffff;
assign target_only_stripe[4323] = 24'hffffff;
assign target_only_stripe[4324] = 24'hffffff;
assign target_only_stripe[4325] = 24'hffffff;
assign target_only_stripe[4326] = 24'hffffff;
assign target_only_stripe[4327] = 24'hffffff;
assign target_only_stripe[4328] = 24'hffffff;
assign target_only_stripe[4329] = 24'hffffff;
assign target_only_stripe[4330] = 24'hffffff;
assign target_only_stripe[4331] = 24'hffffff;
assign target_only_stripe[4332] = 24'hffffff;
assign target_only_stripe[4333] = 24'hffffff;
assign target_only_stripe[4334] = 24'hffffff;
assign target_only_stripe[4335] = 24'hffffff;
assign target_only_stripe[4336] = 24'hffffff;
assign target_only_stripe[4337] = 24'hffffff;
assign target_only_stripe[4338] = 24'hffffff;
assign target_only_stripe[4339] = 24'hffffff;
assign target_only_stripe[4340] = 24'hffffff;
assign target_only_stripe[4341] = 24'hffffff;
assign target_only_stripe[4342] = 24'ha5a5a5;
assign target_only_stripe[4343] = 24'h000000;
assign target_only_stripe[4344] = 24'h000000;
assign target_only_stripe[4345] = 24'h000000;
assign target_only_stripe[4346] = 24'h000000;
assign target_only_stripe[4347] = 24'h000000;
assign target_only_stripe[4348] = 24'h000000;
assign target_only_stripe[4349] = 24'h000000;
assign target_only_stripe[4350] = 24'h000000;
assign target_only_stripe[4351] = 24'h000000;
assign target_only_stripe[4352] = 24'h000000;
assign target_only_stripe[4353] = 24'h000000;
assign target_only_stripe[4354] = 24'h000000;
assign target_only_stripe[4355] = 24'h000000;
assign target_only_stripe[4356] = 24'h000000;
assign target_only_stripe[4357] = 24'h000000;
assign target_only_stripe[4358] = 24'h000000;
assign target_only_stripe[4359] = 24'h000000;
assign target_only_stripe[4360] = 24'h000000;
assign target_only_stripe[4361] = 24'h000000;
assign target_only_stripe[4362] = 24'h000000;
assign target_only_stripe[4363] = 24'h000000;
assign target_only_stripe[4364] = 24'h000000;
assign target_only_stripe[4365] = 24'h000000;
assign target_only_stripe[4366] = 24'h000000;
assign target_only_stripe[4367] = 24'h000000;
assign target_only_stripe[4368] = 24'h000000;
assign target_only_stripe[4369] = 24'h000000;
assign target_only_stripe[4370] = 24'h000000;
assign target_only_stripe[4371] = 24'h000000;
assign target_only_stripe[4372] = 24'h000000;
assign target_only_stripe[4373] = 24'h000000;
assign target_only_stripe[4374] = 24'h000000;
assign target_only_stripe[4375] = 24'h9a9a9a;
assign target_only_stripe[4376] = 24'hffffff;
assign target_only_stripe[4377] = 24'hffffff;
assign target_only_stripe[4378] = 24'hffffff;
assign target_only_stripe[4379] = 24'hffffff;
assign target_only_stripe[4380] = 24'hffffff;
assign target_only_stripe[4381] = 24'hffffff;
assign target_only_stripe[4382] = 24'hffffff;
assign target_only_stripe[4383] = 24'hffffff;
assign target_only_stripe[4384] = 24'hffffff;
assign target_only_stripe[4385] = 24'hffffff;
assign target_only_stripe[4386] = 24'hffffff;
assign target_only_stripe[4387] = 24'hffffff;
assign target_only_stripe[4388] = 24'hffffff;
assign target_only_stripe[4389] = 24'hffffff;
assign target_only_stripe[4390] = 24'hffffff;
assign target_only_stripe[4391] = 24'hffffff;
assign target_only_stripe[4392] = 24'hffffff;
assign target_only_stripe[4393] = 24'hffffff;
assign target_only_stripe[4394] = 24'hffffff;
assign target_only_stripe[4395] = 24'hffffff;
assign target_only_stripe[4396] = 24'hffffff;
assign target_only_stripe[4397] = 24'hffffff;
assign target_only_stripe[4398] = 24'hffffff;
assign target_only_stripe[4399] = 24'hffffff;
assign target_only_stripe[4400] = 24'hffffff;
assign target_only_stripe[4401] = 24'hffffff;
assign target_only_stripe[4402] = 24'hffffff;
assign target_only_stripe[4403] = 24'hffffff;
assign target_only_stripe[4404] = 24'hffffff;
assign target_only_stripe[4405] = 24'hffffff;
assign target_only_stripe[4406] = 24'hffffff;
assign target_only_stripe[4407] = 24'hffffff;
assign target_only_stripe[4408] = 24'hffffff;
assign target_only_stripe[4409] = 24'h4a4a4a;
assign target_only_stripe[4410] = 24'h000000;
assign target_only_stripe[4411] = 24'h000000;
assign target_only_stripe[4412] = 24'h000000;
assign target_only_stripe[4413] = 24'h000000;
assign target_only_stripe[4414] = 24'h000000;
assign target_only_stripe[4415] = 24'h000000;
assign target_only_stripe[4416] = 24'h000000;
assign target_only_stripe[4417] = 24'h000000;
assign target_only_stripe[4418] = 24'h000000;
assign target_only_stripe[4419] = 24'h000000;
assign target_only_stripe[4420] = 24'h000000;
assign target_only_stripe[4421] = 24'h000000;
assign target_only_stripe[4422] = 24'h000000;
assign target_only_stripe[4423] = 24'h000000;
assign target_only_stripe[4424] = 24'h000000;
assign target_only_stripe[4425] = 24'h000000;
assign target_only_stripe[4426] = 24'h000000;
assign target_only_stripe[4427] = 24'h000000;
assign target_only_stripe[4428] = 24'h000000;
assign target_only_stripe[4429] = 24'h000000;
assign target_only_stripe[4430] = 24'h000000;
assign target_only_stripe[4431] = 24'h000000;
assign target_only_stripe[4432] = 24'h000000;
assign target_only_stripe[4433] = 24'h000000;
assign target_only_stripe[4434] = 24'h000000;
assign target_only_stripe[4435] = 24'h000000;
assign target_only_stripe[4436] = 24'h000000;
assign target_only_stripe[4437] = 24'h000000;
assign target_only_stripe[4438] = 24'h000000;
assign target_only_stripe[4439] = 24'h000000;
assign target_only_stripe[4440] = 24'h000000;
assign target_only_stripe[4441] = 24'h000000;
assign target_only_stripe[4442] = 24'h000000;
assign target_only_stripe[4443] = 24'h000000;
assign target_only_stripe[4444] = 24'h000000;
assign target_only_stripe[4445] = 24'h000000;
assign target_only_stripe[4446] = 24'h000000;
assign target_only_stripe[4447] = 24'h000000;
assign target_only_stripe[4448] = 24'h000000;
assign target_only_stripe[4449] = 24'h000000;
assign target_only_stripe[4450] = 24'h000000;
assign target_only_stripe[4451] = 24'h000000;
assign target_only_stripe[4452] = 24'h000000;
assign target_only_stripe[4453] = 24'h000000;
assign target_only_stripe[4454] = 24'h000000;
assign target_only_stripe[4455] = 24'h000000;
assign target_only_stripe[4456] = 24'h000000;
assign target_only_stripe[4457] = 24'h000000;
assign target_only_stripe[4458] = 24'h000000;
assign target_only_stripe[4459] = 24'h000000;
assign target_only_stripe[4460] = 24'h000000;
assign target_only_stripe[4461] = 24'h000000;
assign target_only_stripe[4462] = 24'h000000;
assign target_only_stripe[4463] = 24'h000000;
assign target_only_stripe[4464] = 24'h000000;
assign target_only_stripe[4465] = 24'h000000;
assign target_only_stripe[4466] = 24'h000000;
assign target_only_stripe[4467] = 24'h000000;
assign target_only_stripe[4468] = 24'h000000;
assign target_only_stripe[4469] = 24'h000000;
assign target_only_stripe[4470] = 24'h000000;
assign target_only_stripe[4471] = 24'h000000;
assign target_only_stripe[4472] = 24'h000000;
assign target_only_stripe[4473] = 24'h414141;
assign target_only_stripe[4474] = 24'hffffff;
assign target_only_stripe[4475] = 24'hffffff;
assign target_only_stripe[4476] = 24'hffffff;
assign target_only_stripe[4477] = 24'hffffff;
assign target_only_stripe[4478] = 24'hffffff;
assign target_only_stripe[4479] = 24'hffffff;
assign target_only_stripe[4480] = 24'hffffff;
assign target_only_stripe[4481] = 24'hffffff;
assign target_only_stripe[4482] = 24'hffffff;
assign target_only_stripe[4483] = 24'hffffff;
assign target_only_stripe[4484] = 24'hffffff;
assign target_only_stripe[4485] = 24'hffffff;
assign target_only_stripe[4486] = 24'hffffff;
assign target_only_stripe[4487] = 24'hffffff;
assign target_only_stripe[4488] = 24'hffffff;
assign target_only_stripe[4489] = 24'hffffff;
assign target_only_stripe[4490] = 24'hffffff;
assign target_only_stripe[4491] = 24'hffffff;
assign target_only_stripe[4492] = 24'hffffff;
assign target_only_stripe[4493] = 24'hffffff;
assign target_only_stripe[4494] = 24'hffffff;
assign target_only_stripe[4495] = 24'hffffff;
assign target_only_stripe[4496] = 24'hffffff;
assign target_only_stripe[4497] = 24'hffffff;
assign target_only_stripe[4498] = 24'hffffff;
assign target_only_stripe[4499] = 24'hffffff;
assign target_only_stripe[4500] = 24'hffffff;
assign target_only_stripe[4501] = 24'hffffff;
assign target_only_stripe[4502] = 24'hffffff;
assign target_only_stripe[4503] = 24'hffffff;
assign target_only_stripe[4504] = 24'hffffff;
assign target_only_stripe[4505] = 24'hffffff;
assign target_only_stripe[4506] = 24'hffffff;
assign target_only_stripe[4507] = 24'ha1a1a1;
assign target_only_stripe[4508] = 24'h000000;
assign target_only_stripe[4509] = 24'h000000;
assign target_only_stripe[4510] = 24'h000000;
assign target_only_stripe[4511] = 24'h000000;
assign target_only_stripe[4512] = 24'h000000;
assign target_only_stripe[4513] = 24'h000000;
assign target_only_stripe[4514] = 24'h000000;
assign target_only_stripe[4515] = 24'h000000;
assign target_only_stripe[4516] = 24'h000000;
assign target_only_stripe[4517] = 24'h000000;
assign target_only_stripe[4518] = 24'h000000;
assign target_only_stripe[4519] = 24'h000000;
assign target_only_stripe[4520] = 24'h000000;
assign target_only_stripe[4521] = 24'h000000;
assign target_only_stripe[4522] = 24'h000000;
assign target_only_stripe[4523] = 24'h000000;
assign target_only_stripe[4524] = 24'h000000;
assign target_only_stripe[4525] = 24'h000000;
assign target_only_stripe[4526] = 24'h000000;
assign target_only_stripe[4527] = 24'h000000;
assign target_only_stripe[4528] = 24'h000000;
assign target_only_stripe[4529] = 24'h000000;
assign target_only_stripe[4530] = 24'h000000;
assign target_only_stripe[4531] = 24'h000000;
assign target_only_stripe[4532] = 24'h000000;
assign target_only_stripe[4533] = 24'h000000;
assign target_only_stripe[4534] = 24'h000000;
assign target_only_stripe[4535] = 24'h000000;
assign target_only_stripe[4536] = 24'h000000;
assign target_only_stripe[4537] = 24'h000000;
assign target_only_stripe[4538] = 24'h000000;
assign target_only_stripe[4539] = 24'h000000;
assign target_only_stripe[4540] = 24'hbbbbbb;
assign target_only_stripe[4541] = 24'hffffff;
assign target_only_stripe[4542] = 24'hffffff;
assign target_only_stripe[4543] = 24'hffffff;
assign target_only_stripe[4544] = 24'hffffff;
assign target_only_stripe[4545] = 24'hffffff;
assign target_only_stripe[4546] = 24'hffffff;
assign target_only_stripe[4547] = 24'hffffff;
assign target_only_stripe[4548] = 24'hffffff;
assign target_only_stripe[4549] = 24'hffffff;
assign target_only_stripe[4550] = 24'hffffff;
assign target_only_stripe[4551] = 24'hffffff;
assign target_only_stripe[4552] = 24'hffffff;
assign target_only_stripe[4553] = 24'hffffff;
assign target_only_stripe[4554] = 24'hffffff;
assign target_only_stripe[4555] = 24'hffffff;
assign target_only_stripe[4556] = 24'hffffff;
assign target_only_stripe[4557] = 24'hffffff;
assign target_only_stripe[4558] = 24'hffffff;
assign target_only_stripe[4559] = 24'hffffff;
assign target_only_stripe[4560] = 24'hffffff;
assign target_only_stripe[4561] = 24'hffffff;
assign target_only_stripe[4562] = 24'hffffff;
assign target_only_stripe[4563] = 24'hffffff;
assign target_only_stripe[4564] = 24'hffffff;
assign target_only_stripe[4565] = 24'hffffff;
assign target_only_stripe[4566] = 24'hffffff;
assign target_only_stripe[4567] = 24'hffffff;
assign target_only_stripe[4568] = 24'hffffff;
assign target_only_stripe[4569] = 24'hffffff;
assign target_only_stripe[4570] = 24'hffffff;
assign target_only_stripe[4571] = 24'hffffff;
assign target_only_stripe[4572] = 24'hffffff;
assign target_only_stripe[4573] = 24'hd5c0b0;
assign target_only_stripe[4574] = 24'h1b1b1b;
assign target_only_stripe[4575] = 24'h000000;
assign target_only_stripe[4576] = 24'h000000;
assign target_only_stripe[4577] = 24'h000000;
assign target_only_stripe[4578] = 24'h000000;
assign target_only_stripe[4579] = 24'h000000;
assign target_only_stripe[4580] = 24'h000000;
assign target_only_stripe[4581] = 24'h000000;
assign target_only_stripe[4582] = 24'h000000;
assign target_only_stripe[4583] = 24'h000000;
assign target_only_stripe[4584] = 24'h000000;
assign target_only_stripe[4585] = 24'h000000;
assign target_only_stripe[4586] = 24'h000000;
assign target_only_stripe[4587] = 24'h000000;
assign target_only_stripe[4588] = 24'h000000;
assign target_only_stripe[4589] = 24'h000000;
assign target_only_stripe[4590] = 24'h000000;
assign target_only_stripe[4591] = 24'h000000;
assign target_only_stripe[4592] = 24'h000000;
assign target_only_stripe[4593] = 24'h000000;
assign target_only_stripe[4594] = 24'h000000;
assign target_only_stripe[4595] = 24'h000000;
assign target_only_stripe[4596] = 24'h000000;
assign target_only_stripe[4597] = 24'h000000;
assign target_only_stripe[4598] = 24'h000000;
assign target_only_stripe[4599] = 24'h000000;
assign target_only_stripe[4600] = 24'h000000;
assign target_only_stripe[4601] = 24'h000000;
assign target_only_stripe[4602] = 24'h000000;
assign target_only_stripe[4603] = 24'h000000;
assign target_only_stripe[4604] = 24'h000000;
assign target_only_stripe[4605] = 24'h000000;
assign target_only_stripe[4606] = 24'h000000;
assign target_only_stripe[4607] = 24'h000000;
assign target_only_stripe[4608] = 24'h000000;
assign target_only_stripe[4609] = 24'h000000;
assign target_only_stripe[4610] = 24'h000000;
assign target_only_stripe[4611] = 24'h000000;
assign target_only_stripe[4612] = 24'h000000;
assign target_only_stripe[4613] = 24'h000000;
assign target_only_stripe[4614] = 24'h000000;
assign target_only_stripe[4615] = 24'h000000;
assign target_only_stripe[4616] = 24'h000000;
assign target_only_stripe[4617] = 24'h000000;
assign target_only_stripe[4618] = 24'h000000;
assign target_only_stripe[4619] = 24'h000000;
assign target_only_stripe[4620] = 24'h000000;
assign target_only_stripe[4621] = 24'h000000;
assign target_only_stripe[4622] = 24'h000000;
assign target_only_stripe[4623] = 24'h000000;
assign target_only_stripe[4624] = 24'h000000;
assign target_only_stripe[4625] = 24'h000000;
assign target_only_stripe[4626] = 24'h000000;
assign target_only_stripe[4627] = 24'h000000;
assign target_only_stripe[4628] = 24'h000000;
assign target_only_stripe[4629] = 24'h000000;
assign target_only_stripe[4630] = 24'h000000;
assign target_only_stripe[4631] = 24'h000000;
assign target_only_stripe[4632] = 24'h000000;
assign target_only_stripe[4633] = 24'h000000;
assign target_only_stripe[4634] = 24'h000000;
assign target_only_stripe[4635] = 24'h000000;
assign target_only_stripe[4636] = 24'h000000;
assign target_only_stripe[4637] = 24'h121212;
assign target_only_stripe[4638] = 24'he8e6e6;
assign target_only_stripe[4639] = 24'hffffff;
assign target_only_stripe[4640] = 24'hffffff;
assign target_only_stripe[4641] = 24'hffffff;
assign target_only_stripe[4642] = 24'hffffff;
assign target_only_stripe[4643] = 24'hffffff;
assign target_only_stripe[4644] = 24'hffffff;
assign target_only_stripe[4645] = 24'hffffff;
assign target_only_stripe[4646] = 24'hffffff;
assign target_only_stripe[4647] = 24'hffffff;
assign target_only_stripe[4648] = 24'hffffff;
assign target_only_stripe[4649] = 24'hffffff;
assign target_only_stripe[4650] = 24'hffffff;
assign target_only_stripe[4651] = 24'hffffff;
assign target_only_stripe[4652] = 24'hffffff;
assign target_only_stripe[4653] = 24'hffffff;
assign target_only_stripe[4654] = 24'hffffff;
assign target_only_stripe[4655] = 24'hffffff;
assign target_only_stripe[4656] = 24'hffffff;
assign target_only_stripe[4657] = 24'hffffff;
assign target_only_stripe[4658] = 24'hffffff;
assign target_only_stripe[4659] = 24'hffffff;
assign target_only_stripe[4660] = 24'hffffff;
assign target_only_stripe[4661] = 24'hffffff;
assign target_only_stripe[4662] = 24'hffffff;
assign target_only_stripe[4663] = 24'hffffff;
assign target_only_stripe[4664] = 24'hffffff;
assign target_only_stripe[4665] = 24'hffffff;
assign target_only_stripe[4666] = 24'hffffff;
assign target_only_stripe[4667] = 24'hffffff;
assign target_only_stripe[4668] = 24'hffffff;
assign target_only_stripe[4669] = 24'hffffff;
assign target_only_stripe[4670] = 24'hffffff;
assign target_only_stripe[4671] = 24'ha8a8a8;
assign target_only_stripe[4672] = 24'h000000;
assign target_only_stripe[4673] = 24'h000000;
assign target_only_stripe[4674] = 24'h000000;
assign target_only_stripe[4675] = 24'h000000;
assign target_only_stripe[4676] = 24'h000000;
assign target_only_stripe[4677] = 24'h000000;
assign target_only_stripe[4678] = 24'h000000;
assign target_only_stripe[4679] = 24'h000000;
assign target_only_stripe[4680] = 24'h000000;
assign target_only_stripe[4681] = 24'h000000;
assign target_only_stripe[4682] = 24'h000000;
assign target_only_stripe[4683] = 24'h000000;
assign target_only_stripe[4684] = 24'h000000;
assign target_only_stripe[4685] = 24'h000000;
assign target_only_stripe[4686] = 24'h000000;
assign target_only_stripe[4687] = 24'h000000;
assign target_only_stripe[4688] = 24'h000000;
assign target_only_stripe[4689] = 24'h000000;
assign target_only_stripe[4690] = 24'h000000;
assign target_only_stripe[4691] = 24'h000000;
assign target_only_stripe[4692] = 24'h000000;
assign target_only_stripe[4693] = 24'h000000;
assign target_only_stripe[4694] = 24'h000000;
assign target_only_stripe[4695] = 24'h000000;
assign target_only_stripe[4696] = 24'h000000;
assign target_only_stripe[4697] = 24'h000000;
assign target_only_stripe[4698] = 24'h000000;
assign target_only_stripe[4699] = 24'h000000;
assign target_only_stripe[4700] = 24'h000000;
assign target_only_stripe[4701] = 24'h000000;
assign target_only_stripe[4702] = 24'h000000;
assign target_only_stripe[4703] = 24'h000000;
assign target_only_stripe[4704] = 24'h959595;
assign target_only_stripe[4705] = 24'hffffff;
assign target_only_stripe[4706] = 24'hffffff;
assign target_only_stripe[4707] = 24'hffffff;
assign target_only_stripe[4708] = 24'hffffff;
assign target_only_stripe[4709] = 24'hffffff;
assign target_only_stripe[4710] = 24'hffffff;
assign target_only_stripe[4711] = 24'hffffff;
assign target_only_stripe[4712] = 24'hffffff;
assign target_only_stripe[4713] = 24'hffffff;
assign target_only_stripe[4714] = 24'hffffff;
assign target_only_stripe[4715] = 24'hffffff;
assign target_only_stripe[4716] = 24'hffffff;
assign target_only_stripe[4717] = 24'hffffff;
assign target_only_stripe[4718] = 24'hffffff;
assign target_only_stripe[4719] = 24'hffffff;
assign target_only_stripe[4720] = 24'hffffff;
assign target_only_stripe[4721] = 24'hffffff;
assign target_only_stripe[4722] = 24'hffffff;
assign target_only_stripe[4723] = 24'hffffff;
assign target_only_stripe[4724] = 24'hffffff;
assign target_only_stripe[4725] = 24'hffffff;
assign target_only_stripe[4726] = 24'hffffff;
assign target_only_stripe[4727] = 24'hffffff;
assign target_only_stripe[4728] = 24'hffffff;
assign target_only_stripe[4729] = 24'hffffff;
assign target_only_stripe[4730] = 24'hffffff;
assign target_only_stripe[4731] = 24'hffffff;
assign target_only_stripe[4732] = 24'hffffff;
assign target_only_stripe[4733] = 24'hffffff;
assign target_only_stripe[4734] = 24'hffffff;
assign target_only_stripe[4735] = 24'hffffff;
assign target_only_stripe[4736] = 24'hffffff;
assign target_only_stripe[4737] = 24'hffffff;
assign target_only_stripe[4738] = 24'hffffff;
assign target_only_stripe[4739] = 24'h000000;
assign target_only_stripe[4740] = 24'h000000;
assign target_only_stripe[4741] = 24'h000000;
assign target_only_stripe[4742] = 24'h000000;
assign target_only_stripe[4743] = 24'h000000;
assign target_only_stripe[4744] = 24'h000000;
assign target_only_stripe[4745] = 24'h000000;
assign target_only_stripe[4746] = 24'h000000;
assign target_only_stripe[4747] = 24'h000000;
assign target_only_stripe[4748] = 24'h000000;
assign target_only_stripe[4749] = 24'h000000;
assign target_only_stripe[4750] = 24'h000000;
assign target_only_stripe[4751] = 24'h000000;
assign target_only_stripe[4752] = 24'h000000;
assign target_only_stripe[4753] = 24'h000000;
assign target_only_stripe[4754] = 24'h000000;
assign target_only_stripe[4755] = 24'h000000;
assign target_only_stripe[4756] = 24'h000000;
assign target_only_stripe[4757] = 24'h000000;
assign target_only_stripe[4758] = 24'h000000;
assign target_only_stripe[4759] = 24'h000000;
assign target_only_stripe[4760] = 24'h000000;
assign target_only_stripe[4761] = 24'h000000;
assign target_only_stripe[4762] = 24'h000000;
assign target_only_stripe[4763] = 24'h000000;
assign target_only_stripe[4764] = 24'h000000;
assign target_only_stripe[4765] = 24'h000000;
assign target_only_stripe[4766] = 24'h000000;
assign target_only_stripe[4767] = 24'h000000;
assign target_only_stripe[4768] = 24'h000000;
assign target_only_stripe[4769] = 24'h000000;
assign target_only_stripe[4770] = 24'h000000;
assign target_only_stripe[4771] = 24'h000000;
assign target_only_stripe[4772] = 24'h000000;
assign target_only_stripe[4773] = 24'h000000;
assign target_only_stripe[4774] = 24'h000000;
assign target_only_stripe[4775] = 24'h000000;
assign target_only_stripe[4776] = 24'h000000;
assign target_only_stripe[4777] = 24'h000000;
assign target_only_stripe[4778] = 24'h000000;
assign target_only_stripe[4779] = 24'h000000;
assign target_only_stripe[4780] = 24'h000000;
assign target_only_stripe[4781] = 24'h000000;
assign target_only_stripe[4782] = 24'h000000;
assign target_only_stripe[4783] = 24'h000000;
assign target_only_stripe[4784] = 24'h000000;
assign target_only_stripe[4785] = 24'h000000;
assign target_only_stripe[4786] = 24'h000000;
assign target_only_stripe[4787] = 24'h000000;
assign target_only_stripe[4788] = 24'h000000;
assign target_only_stripe[4789] = 24'h000000;
assign target_only_stripe[4790] = 24'h000000;
assign target_only_stripe[4791] = 24'h000000;
assign target_only_stripe[4792] = 24'h000000;
assign target_only_stripe[4793] = 24'h000000;
assign target_only_stripe[4794] = 24'h000000;
assign target_only_stripe[4795] = 24'h000000;
assign target_only_stripe[4796] = 24'h000000;
assign target_only_stripe[4797] = 24'h000000;
assign target_only_stripe[4798] = 24'h000000;
assign target_only_stripe[4799] = 24'h000000;
assign target_only_stripe[4800] = 24'h000000;
assign target_only_stripe[4801] = 24'h000000;
assign target_only_stripe[4802] = 24'hffffff;
assign target_only_stripe[4803] = 24'hffffff;
assign target_only_stripe[4804] = 24'hffffff;
assign target_only_stripe[4805] = 24'hffffff;
assign target_only_stripe[4806] = 24'hffffff;
assign target_only_stripe[4807] = 24'hffffff;
assign target_only_stripe[4808] = 24'hffffff;
assign target_only_stripe[4809] = 24'hffffff;
assign target_only_stripe[4810] = 24'hffffff;
assign target_only_stripe[4811] = 24'hffffff;
assign target_only_stripe[4812] = 24'hffffff;
assign target_only_stripe[4813] = 24'hffffff;
assign target_only_stripe[4814] = 24'hffffff;
assign target_only_stripe[4815] = 24'hffffff;
assign target_only_stripe[4816] = 24'hffffff;
assign target_only_stripe[4817] = 24'hffffff;
assign target_only_stripe[4818] = 24'hffffff;
assign target_only_stripe[4819] = 24'hffffff;
assign target_only_stripe[4820] = 24'hffffff;
assign target_only_stripe[4821] = 24'hffffff;
assign target_only_stripe[4822] = 24'hffffff;
assign target_only_stripe[4823] = 24'hffffff;
assign target_only_stripe[4824] = 24'hffffff;
assign target_only_stripe[4825] = 24'hffffff;
assign target_only_stripe[4826] = 24'hffffff;
assign target_only_stripe[4827] = 24'hffffff;
assign target_only_stripe[4828] = 24'hffffff;
assign target_only_stripe[4829] = 24'hffffff;
assign target_only_stripe[4830] = 24'hffffff;
assign target_only_stripe[4831] = 24'hffffff;
assign target_only_stripe[4832] = 24'hffffff;
assign target_only_stripe[4833] = 24'hffffff;
assign target_only_stripe[4834] = 24'hffffff;
assign target_only_stripe[4835] = 24'hffffff;
assign target_only_stripe[4836] = 24'h9d9d9d;
assign target_only_stripe[4837] = 24'h000000;
assign target_only_stripe[4838] = 24'h000000;
assign target_only_stripe[4839] = 24'h000000;
assign target_only_stripe[4840] = 24'h000000;
assign target_only_stripe[4841] = 24'h000000;
assign target_only_stripe[4842] = 24'h000000;
assign target_only_stripe[4843] = 24'h000000;
assign target_only_stripe[4844] = 24'h000000;
assign target_only_stripe[4845] = 24'h000000;
assign target_only_stripe[4846] = 24'h000000;
assign target_only_stripe[4847] = 24'h000000;
assign target_only_stripe[4848] = 24'h000000;
assign target_only_stripe[4849] = 24'h000000;
assign target_only_stripe[4850] = 24'h000000;
assign target_only_stripe[4851] = 24'h000000;
assign target_only_stripe[4852] = 24'h000000;
assign target_only_stripe[4853] = 24'h000000;
assign target_only_stripe[4854] = 24'h000000;
assign target_only_stripe[4855] = 24'h000000;
assign target_only_stripe[4856] = 24'h000000;
assign target_only_stripe[4857] = 24'h000000;
assign target_only_stripe[4858] = 24'h000000;
assign target_only_stripe[4859] = 24'h000000;
assign target_only_stripe[4860] = 24'h000000;
assign target_only_stripe[4861] = 24'h000000;
assign target_only_stripe[4862] = 24'h000000;
assign target_only_stripe[4863] = 24'h000000;
assign target_only_stripe[4864] = 24'h000000;
assign target_only_stripe[4865] = 24'h000000;
assign target_only_stripe[4866] = 24'h000000;
assign target_only_stripe[4867] = 24'h000000;
assign target_only_stripe[4868] = 24'h000000;
assign target_only_stripe[4869] = 24'ha1a1a1;
assign target_only_stripe[4870] = 24'hffffff;
assign target_only_stripe[4871] = 24'hffffff;
assign target_only_stripe[4872] = 24'hffffff;
assign target_only_stripe[4873] = 24'hffffff;
assign target_only_stripe[4874] = 24'hffffff;
assign target_only_stripe[4875] = 24'hffffff;
assign target_only_stripe[4876] = 24'hffffff;
assign target_only_stripe[4877] = 24'hffffff;
assign target_only_stripe[4878] = 24'hffffff;
assign target_only_stripe[4879] = 24'hffffff;
assign target_only_stripe[4880] = 24'hffffff;
assign target_only_stripe[4881] = 24'hffffff;
assign target_only_stripe[4882] = 24'hffffff;
assign target_only_stripe[4883] = 24'hffffff;
assign target_only_stripe[4884] = 24'hffffff;
assign target_only_stripe[4885] = 24'hffffff;
assign target_only_stripe[4886] = 24'hffffff;
assign target_only_stripe[4887] = 24'hffffff;
assign target_only_stripe[4888] = 24'hffffff;
assign target_only_stripe[4889] = 24'hffffff;
assign target_only_stripe[4890] = 24'hffffff;
assign target_only_stripe[4891] = 24'hffffff;
assign target_only_stripe[4892] = 24'hffffff;
assign target_only_stripe[4893] = 24'hffffff;
assign target_only_stripe[4894] = 24'hffffff;
assign target_only_stripe[4895] = 24'hffffff;
assign target_only_stripe[4896] = 24'hffffff;
assign target_only_stripe[4897] = 24'hffffff;
assign target_only_stripe[4898] = 24'hffffff;
assign target_only_stripe[4899] = 24'hffffff;
assign target_only_stripe[4900] = 24'hffffff;
assign target_only_stripe[4901] = 24'hffffff;
assign target_only_stripe[4902] = 24'hddc6b3;
assign target_only_stripe[4903] = 24'h1b1b1b;
assign target_only_stripe[4904] = 24'h000000;
assign target_only_stripe[4905] = 24'h000000;
assign target_only_stripe[4906] = 24'h000000;
assign target_only_stripe[4907] = 24'h000000;
assign target_only_stripe[4908] = 24'h000000;
assign target_only_stripe[4909] = 24'h000000;
assign target_only_stripe[4910] = 24'h000000;
assign target_only_stripe[4911] = 24'h000000;
assign target_only_stripe[4912] = 24'h000000;
assign target_only_stripe[4913] = 24'h000000;
assign target_only_stripe[4914] = 24'h000000;
assign target_only_stripe[4915] = 24'h000000;
assign target_only_stripe[4916] = 24'h000000;
assign target_only_stripe[4917] = 24'h000000;
assign target_only_stripe[4918] = 24'h000000;
assign target_only_stripe[4919] = 24'h000000;
assign target_only_stripe[4920] = 24'h000000;
assign target_only_stripe[4921] = 24'h000000;
assign target_only_stripe[4922] = 24'h000000;
assign target_only_stripe[4923] = 24'h000000;
assign target_only_stripe[4924] = 24'h000000;
assign target_only_stripe[4925] = 24'h000000;
assign target_only_stripe[4926] = 24'h000000;
assign target_only_stripe[4927] = 24'h000000;
assign target_only_stripe[4928] = 24'h000000;
assign target_only_stripe[4929] = 24'h000000;
assign target_only_stripe[4930] = 24'h000000;
assign target_only_stripe[4931] = 24'h000000;
assign target_only_stripe[4932] = 24'h000000;
assign target_only_stripe[4933] = 24'h000000;
assign target_only_stripe[4934] = 24'h000000;
assign target_only_stripe[4935] = 24'h000000;
assign target_only_stripe[4936] = 24'h000000;
assign target_only_stripe[4937] = 24'h000000;
assign target_only_stripe[4938] = 24'h000000;
assign target_only_stripe[4939] = 24'h000000;
assign target_only_stripe[4940] = 24'h000000;
assign target_only_stripe[4941] = 24'h000000;
assign target_only_stripe[4942] = 24'h000000;
assign target_only_stripe[4943] = 24'h000000;
assign target_only_stripe[4944] = 24'h000000;
assign target_only_stripe[4945] = 24'h000000;
assign target_only_stripe[4946] = 24'h000000;
assign target_only_stripe[4947] = 24'h000000;
assign target_only_stripe[4948] = 24'h000000;
assign target_only_stripe[4949] = 24'h000000;
assign target_only_stripe[4950] = 24'h000000;
assign target_only_stripe[4951] = 24'h000000;
assign target_only_stripe[4952] = 24'h000000;
assign target_only_stripe[4953] = 24'h000000;
assign target_only_stripe[4954] = 24'h000000;
assign target_only_stripe[4955] = 24'h000000;
assign target_only_stripe[4956] = 24'h000000;
assign target_only_stripe[4957] = 24'h000000;
assign target_only_stripe[4958] = 24'h000000;
assign target_only_stripe[4959] = 24'h000000;
assign target_only_stripe[4960] = 24'h000000;
assign target_only_stripe[4961] = 24'h000000;
assign target_only_stripe[4962] = 24'h000000;
assign target_only_stripe[4963] = 24'h000000;
assign target_only_stripe[4964] = 24'h000000;
assign target_only_stripe[4965] = 24'h000000;
assign target_only_stripe[4966] = 24'h111111;
assign target_only_stripe[4967] = 24'he9e9e9;
assign target_only_stripe[4968] = 24'hffffff;
assign target_only_stripe[4969] = 24'hffffff;
assign target_only_stripe[4970] = 24'hffffff;
assign target_only_stripe[4971] = 24'hffffff;
assign target_only_stripe[4972] = 24'hffffff;
assign target_only_stripe[4973] = 24'hffffff;
assign target_only_stripe[4974] = 24'hffffff;
assign target_only_stripe[4975] = 24'hffffff;
assign target_only_stripe[4976] = 24'hffffff;
assign target_only_stripe[4977] = 24'hffffff;
assign target_only_stripe[4978] = 24'hffffff;
assign target_only_stripe[4979] = 24'hffffff;
assign target_only_stripe[4980] = 24'hffffff;
assign target_only_stripe[4981] = 24'hffffff;
assign target_only_stripe[4982] = 24'hffffff;
assign target_only_stripe[4983] = 24'hffffff;
assign target_only_stripe[4984] = 24'hffffff;
assign target_only_stripe[4985] = 24'hffffff;
assign target_only_stripe[4986] = 24'hffffff;
assign target_only_stripe[4987] = 24'hffffff;
assign target_only_stripe[4988] = 24'hffffff;
assign target_only_stripe[4989] = 24'hffffff;
assign target_only_stripe[4990] = 24'hffffff;
assign target_only_stripe[4991] = 24'hffffff;
assign target_only_stripe[4992] = 24'hffffff;
assign target_only_stripe[4993] = 24'hffffff;
assign target_only_stripe[4994] = 24'hffffff;
assign target_only_stripe[4995] = 24'hffffff;
assign target_only_stripe[4996] = 24'hffffff;
assign target_only_stripe[4997] = 24'hffffff;
assign target_only_stripe[4998] = 24'hffffff;
assign target_only_stripe[4999] = 24'hffffff;
assign target_only_stripe[5000] = 24'hbbbbbb;
assign target_only_stripe[5001] = 24'h000000;
assign target_only_stripe[5002] = 24'h000000;
assign target_only_stripe[5003] = 24'h000000;
assign target_only_stripe[5004] = 24'h000000;
assign target_only_stripe[5005] = 24'h000000;
assign target_only_stripe[5006] = 24'h000000;
assign target_only_stripe[5007] = 24'h000000;
assign target_only_stripe[5008] = 24'h000000;
assign target_only_stripe[5009] = 24'h000000;
assign target_only_stripe[5010] = 24'h000000;
assign target_only_stripe[5011] = 24'h000000;
assign target_only_stripe[5012] = 24'h000000;
assign target_only_stripe[5013] = 24'h000000;
assign target_only_stripe[5014] = 24'h000000;
assign target_only_stripe[5015] = 24'h000000;
assign target_only_stripe[5016] = 24'h000000;
assign target_only_stripe[5017] = 24'h000000;
assign target_only_stripe[5018] = 24'h000000;
assign target_only_stripe[5019] = 24'h000000;
assign target_only_stripe[5020] = 24'h000000;
assign target_only_stripe[5021] = 24'h000000;
assign target_only_stripe[5022] = 24'h000000;
assign target_only_stripe[5023] = 24'h000000;
assign target_only_stripe[5024] = 24'h000000;
assign target_only_stripe[5025] = 24'h000000;
assign target_only_stripe[5026] = 24'h000000;
assign target_only_stripe[5027] = 24'h000000;
assign target_only_stripe[5028] = 24'h000000;
assign target_only_stripe[5029] = 24'h000000;
assign target_only_stripe[5030] = 24'h000000;
assign target_only_stripe[5031] = 24'h000000;
assign target_only_stripe[5032] = 24'h000000;
assign target_only_stripe[5033] = 24'h8b8b8b;
assign target_only_stripe[5034] = 24'hffffff;
assign target_only_stripe[5035] = 24'hffffff;
assign target_only_stripe[5036] = 24'hffffff;
assign target_only_stripe[5037] = 24'hffffff;
assign target_only_stripe[5038] = 24'hffffff;
assign target_only_stripe[5039] = 24'hffffff;
assign target_only_stripe[5040] = 24'hffffff;
assign target_only_stripe[5041] = 24'hffffff;
assign target_only_stripe[5042] = 24'hffffff;
assign target_only_stripe[5043] = 24'hffffff;
assign target_only_stripe[5044] = 24'hffffff;
assign target_only_stripe[5045] = 24'hffffff;
assign target_only_stripe[5046] = 24'hffffff;
assign target_only_stripe[5047] = 24'hffffff;
assign target_only_stripe[5048] = 24'hffffff;
assign target_only_stripe[5049] = 24'hffffff;
assign target_only_stripe[5050] = 24'hffffff;
assign target_only_stripe[5051] = 24'hffffff;
assign target_only_stripe[5052] = 24'hffffff;
assign target_only_stripe[5053] = 24'hffffff;
assign target_only_stripe[5054] = 24'hffffff;
assign target_only_stripe[5055] = 24'hffffff;
assign target_only_stripe[5056] = 24'hffffff;
assign target_only_stripe[5057] = 24'hffffff;
assign target_only_stripe[5058] = 24'hffffff;
assign target_only_stripe[5059] = 24'hffffff;
assign target_only_stripe[5060] = 24'hffffff;
assign target_only_stripe[5061] = 24'hffffff;
assign target_only_stripe[5062] = 24'hffffff;
assign target_only_stripe[5063] = 24'hffffff;
assign target_only_stripe[5064] = 24'hffffff;
assign target_only_stripe[5065] = 24'hffffff;
assign target_only_stripe[5066] = 24'hffffff;
assign target_only_stripe[5067] = 24'hffffff;
assign target_only_stripe[5068] = 24'h000000;
assign target_only_stripe[5069] = 24'h000000;
assign target_only_stripe[5070] = 24'h000000;
assign target_only_stripe[5071] = 24'h000000;
assign target_only_stripe[5072] = 24'h000000;
assign target_only_stripe[5073] = 24'h000000;
assign target_only_stripe[5074] = 24'h000000;
assign target_only_stripe[5075] = 24'h000000;
assign target_only_stripe[5076] = 24'h000000;
assign target_only_stripe[5077] = 24'h000000;
assign target_only_stripe[5078] = 24'h000000;
assign target_only_stripe[5079] = 24'h000000;
assign target_only_stripe[5080] = 24'h000000;
assign target_only_stripe[5081] = 24'h000000;
assign target_only_stripe[5082] = 24'h000000;
assign target_only_stripe[5083] = 24'h000000;
assign target_only_stripe[5084] = 24'h000000;
assign target_only_stripe[5085] = 24'h000000;
assign target_only_stripe[5086] = 24'h000000;
assign target_only_stripe[5087] = 24'h000000;
assign target_only_stripe[5088] = 24'h000000;
assign target_only_stripe[5089] = 24'h000000;
assign target_only_stripe[5090] = 24'h000000;
assign target_only_stripe[5091] = 24'h000000;
assign target_only_stripe[5092] = 24'h000000;
assign target_only_stripe[5093] = 24'h000000;
assign target_only_stripe[5094] = 24'h000000;
assign target_only_stripe[5095] = 24'h000000;
assign target_only_stripe[5096] = 24'h000000;
assign target_only_stripe[5097] = 24'h000000;
assign target_only_stripe[5098] = 24'h000000;
assign target_only_stripe[5099] = 24'h000000;
assign target_only_stripe[5100] = 24'h000000;
assign target_only_stripe[5101] = 24'h000000;
assign target_only_stripe[5102] = 24'h000000;
assign target_only_stripe[5103] = 24'h000000;
assign target_only_stripe[5104] = 24'h000000;
assign target_only_stripe[5105] = 24'h000000;
assign target_only_stripe[5106] = 24'h000000;
assign target_only_stripe[5107] = 24'h000000;
assign target_only_stripe[5108] = 24'h000000;
assign target_only_stripe[5109] = 24'h000000;
assign target_only_stripe[5110] = 24'h000000;
assign target_only_stripe[5111] = 24'h000000;
assign target_only_stripe[5112] = 24'h000000;
assign target_only_stripe[5113] = 24'h000000;
assign target_only_stripe[5114] = 24'h000000;
assign target_only_stripe[5115] = 24'h000000;
assign target_only_stripe[5116] = 24'h000000;
assign target_only_stripe[5117] = 24'h000000;
assign target_only_stripe[5118] = 24'h000000;
assign target_only_stripe[5119] = 24'h000000;
assign target_only_stripe[5120] = 24'h000000;
assign target_only_stripe[5121] = 24'h000000;
assign target_only_stripe[5122] = 24'h000000;
assign target_only_stripe[5123] = 24'h000000;
assign target_only_stripe[5124] = 24'h000000;
assign target_only_stripe[5125] = 24'h000000;
assign target_only_stripe[5126] = 24'h000000;
assign target_only_stripe[5127] = 24'h000000;
assign target_only_stripe[5128] = 24'h000000;
assign target_only_stripe[5129] = 24'h000000;
assign target_only_stripe[5130] = 24'h000000;
assign target_only_stripe[5131] = 24'hffffff;
assign target_only_stripe[5132] = 24'hffffff;
assign target_only_stripe[5133] = 24'hffffff;
assign target_only_stripe[5134] = 24'hffffff;
assign target_only_stripe[5135] = 24'hffffff;
assign target_only_stripe[5136] = 24'hffffff;
assign target_only_stripe[5137] = 24'hffffff;
assign target_only_stripe[5138] = 24'hffffff;
assign target_only_stripe[5139] = 24'hffffff;
assign target_only_stripe[5140] = 24'hffffff;
assign target_only_stripe[5141] = 24'hffffff;
assign target_only_stripe[5142] = 24'hffffff;
assign target_only_stripe[5143] = 24'hffffff;
assign target_only_stripe[5144] = 24'hffffff;
assign target_only_stripe[5145] = 24'hffffff;
assign target_only_stripe[5146] = 24'hffffff;
assign target_only_stripe[5147] = 24'hffffff;
assign target_only_stripe[5148] = 24'hffffff;
assign target_only_stripe[5149] = 24'hffffff;
assign target_only_stripe[5150] = 24'hffffff;
assign target_only_stripe[5151] = 24'hffffff;
assign target_only_stripe[5152] = 24'hffffff;
assign target_only_stripe[5153] = 24'hffffff;
assign target_only_stripe[5154] = 24'hffffff;
assign target_only_stripe[5155] = 24'hffffff;
assign target_only_stripe[5156] = 24'hffffff;
assign target_only_stripe[5157] = 24'hffffff;
assign target_only_stripe[5158] = 24'hffffff;
assign target_only_stripe[5159] = 24'hffffff;
assign target_only_stripe[5160] = 24'hffffff;
assign target_only_stripe[5161] = 24'hffffff;
assign target_only_stripe[5162] = 24'hffffff;
assign target_only_stripe[5163] = 24'hffffff;
assign target_only_stripe[5164] = 24'hffffff;
assign target_only_stripe[5165] = 24'h939393;
assign target_only_stripe[5166] = 24'h000000;
assign target_only_stripe[5167] = 24'h000000;
assign target_only_stripe[5168] = 24'h000000;
assign target_only_stripe[5169] = 24'h000000;
assign target_only_stripe[5170] = 24'h000000;
assign target_only_stripe[5171] = 24'h000000;
assign target_only_stripe[5172] = 24'h000000;
assign target_only_stripe[5173] = 24'h000000;
assign target_only_stripe[5174] = 24'h000000;
assign target_only_stripe[5175] = 24'h000000;
assign target_only_stripe[5176] = 24'h000000;
assign target_only_stripe[5177] = 24'h000000;
assign target_only_stripe[5178] = 24'h000000;
assign target_only_stripe[5179] = 24'h000000;
assign target_only_stripe[5180] = 24'h000000;
assign target_only_stripe[5181] = 24'h000000;
assign target_only_stripe[5182] = 24'h000000;
assign target_only_stripe[5183] = 24'h000000;
assign target_only_stripe[5184] = 24'h000000;
assign target_only_stripe[5185] = 24'h000000;
assign target_only_stripe[5186] = 24'h000000;
assign target_only_stripe[5187] = 24'h000000;
assign target_only_stripe[5188] = 24'h000000;
assign target_only_stripe[5189] = 24'h000000;
assign target_only_stripe[5190] = 24'h000000;
assign target_only_stripe[5191] = 24'h000000;
assign target_only_stripe[5192] = 24'h000000;
assign target_only_stripe[5193] = 24'h000000;
assign target_only_stripe[5194] = 24'h000000;
assign target_only_stripe[5195] = 24'h000000;
assign target_only_stripe[5196] = 24'h000000;
assign target_only_stripe[5197] = 24'h000000;
assign target_only_stripe[5198] = 24'hb4b4b4;
assign target_only_stripe[5199] = 24'hffffff;
assign target_only_stripe[5200] = 24'hffffff;
assign target_only_stripe[5201] = 24'hffffff;
assign target_only_stripe[5202] = 24'hffffff;
assign target_only_stripe[5203] = 24'hffffff;
assign target_only_stripe[5204] = 24'hffffff;
assign target_only_stripe[5205] = 24'hffffff;
assign target_only_stripe[5206] = 24'hffffff;
assign target_only_stripe[5207] = 24'hffffff;
assign target_only_stripe[5208] = 24'hffffff;
assign target_only_stripe[5209] = 24'hffffff;
assign target_only_stripe[5210] = 24'hffffff;
assign target_only_stripe[5211] = 24'hffffff;
assign target_only_stripe[5212] = 24'hffffff;
assign target_only_stripe[5213] = 24'hffffff;
assign target_only_stripe[5214] = 24'hffffff;
assign target_only_stripe[5215] = 24'hffffff;
assign target_only_stripe[5216] = 24'hffffff;
assign target_only_stripe[5217] = 24'hffffff;
assign target_only_stripe[5218] = 24'hffffff;
assign target_only_stripe[5219] = 24'hffffff;
assign target_only_stripe[5220] = 24'hffffff;
assign target_only_stripe[5221] = 24'hffffff;
assign target_only_stripe[5222] = 24'hfaf7f5;
assign target_only_stripe[5223] = 24'hffffff;
assign target_only_stripe[5224] = 24'hffffff;
assign target_only_stripe[5225] = 24'hfaf7f5;
assign target_only_stripe[5226] = 24'hffffff;
assign target_only_stripe[5227] = 24'hffffff;
assign target_only_stripe[5228] = 24'hffffff;
assign target_only_stripe[5229] = 24'hffffff;
assign target_only_stripe[5230] = 24'hfaf7f5;
assign target_only_stripe[5231] = 24'hdfd2c8;
assign target_only_stripe[5232] = 24'h1b1b1b;
assign target_only_stripe[5233] = 24'h000000;
assign target_only_stripe[5234] = 24'h000000;
assign target_only_stripe[5235] = 24'h000000;
assign target_only_stripe[5236] = 24'h000000;
assign target_only_stripe[5237] = 24'h000000;
assign target_only_stripe[5238] = 24'h000000;
assign target_only_stripe[5239] = 24'h000000;
assign target_only_stripe[5240] = 24'h000000;
assign target_only_stripe[5241] = 24'h000000;
assign target_only_stripe[5242] = 24'h000000;
assign target_only_stripe[5243] = 24'h000000;
assign target_only_stripe[5244] = 24'h000000;
assign target_only_stripe[5245] = 24'h000000;
assign target_only_stripe[5246] = 24'h000000;
assign target_only_stripe[5247] = 24'h000000;
assign target_only_stripe[5248] = 24'h000000;
assign target_only_stripe[5249] = 24'h000000;
assign target_only_stripe[5250] = 24'h000000;
assign target_only_stripe[5251] = 24'h000000;
assign target_only_stripe[5252] = 24'h000000;
assign target_only_stripe[5253] = 24'h000000;
assign target_only_stripe[5254] = 24'h000000;
assign target_only_stripe[5255] = 24'h000000;
assign target_only_stripe[5256] = 24'h000000;
assign target_only_stripe[5257] = 24'h000000;
assign target_only_stripe[5258] = 24'h000000;
assign target_only_stripe[5259] = 24'h000000;
assign target_only_stripe[5260] = 24'h000000;
assign target_only_stripe[5261] = 24'h000000;
assign target_only_stripe[5262] = 24'h000000;
assign target_only_stripe[5263] = 24'h000000;
assign target_only_stripe[5264] = 24'h000000;
assign target_only_stripe[5265] = 24'h000000;
assign target_only_stripe[5266] = 24'h000000;
assign target_only_stripe[5267] = 24'h000000;
assign target_only_stripe[5268] = 24'h000000;
assign target_only_stripe[5269] = 24'h000000;
assign target_only_stripe[5270] = 24'h000000;
assign target_only_stripe[5271] = 24'h000000;
assign target_only_stripe[5272] = 24'h000000;
assign target_only_stripe[5273] = 24'h000000;
assign target_only_stripe[5274] = 24'h000000;
assign target_only_stripe[5275] = 24'h000000;
assign target_only_stripe[5276] = 24'h000000;
assign target_only_stripe[5277] = 24'h000000;
assign target_only_stripe[5278] = 24'h000000;
assign target_only_stripe[5279] = 24'h000000;
assign target_only_stripe[5280] = 24'h000000;
assign target_only_stripe[5281] = 24'h000000;
assign target_only_stripe[5282] = 24'h000000;
assign target_only_stripe[5283] = 24'h000000;
assign target_only_stripe[5284] = 24'h000000;
assign target_only_stripe[5285] = 24'h000000;
assign target_only_stripe[5286] = 24'h000000;
assign target_only_stripe[5287] = 24'h000000;
assign target_only_stripe[5288] = 24'h000000;
assign target_only_stripe[5289] = 24'h000000;
assign target_only_stripe[5290] = 24'h000000;
assign target_only_stripe[5291] = 24'h000000;
assign target_only_stripe[5292] = 24'h000000;
assign target_only_stripe[5293] = 24'h000000;
assign target_only_stripe[5294] = 24'h000000;
assign target_only_stripe[5295] = 24'h101010;
assign target_only_stripe[5296] = 24'he5e5e5;
assign target_only_stripe[5297] = 24'hffffff;
assign target_only_stripe[5298] = 24'hffffff;
assign target_only_stripe[5299] = 24'hffffff;
assign target_only_stripe[5300] = 24'hffffff;
assign target_only_stripe[5301] = 24'hffffff;
assign target_only_stripe[5302] = 24'hffffff;
assign target_only_stripe[5303] = 24'hffffff;
assign target_only_stripe[5304] = 24'hffffff;
assign target_only_stripe[5305] = 24'hffffff;
assign target_only_stripe[5306] = 24'hffffff;
assign target_only_stripe[5307] = 24'hffffff;
assign target_only_stripe[5308] = 24'hffffff;
assign target_only_stripe[5309] = 24'hffffff;
assign target_only_stripe[5310] = 24'hffffff;
assign target_only_stripe[5311] = 24'hffffff;
assign target_only_stripe[5312] = 24'hffffff;
assign target_only_stripe[5313] = 24'hffffff;
assign target_only_stripe[5314] = 24'hffffff;
assign target_only_stripe[5315] = 24'hffffff;
assign target_only_stripe[5316] = 24'hffffff;
assign target_only_stripe[5317] = 24'hffffff;
assign target_only_stripe[5318] = 24'hffffff;
assign target_only_stripe[5319] = 24'hffffff;
assign target_only_stripe[5320] = 24'hffffff;
assign target_only_stripe[5321] = 24'hffffff;
assign target_only_stripe[5322] = 24'hffffff;
assign target_only_stripe[5323] = 24'hffffff;
assign target_only_stripe[5324] = 24'hffffff;
assign target_only_stripe[5325] = 24'hffffff;
assign target_only_stripe[5326] = 24'hffffff;
assign target_only_stripe[5327] = 24'hffffff;
assign target_only_stripe[5328] = 24'hffffff;
assign target_only_stripe[5329] = 24'hc9c9c9;
assign target_only_stripe[5330] = 24'h000000;
assign target_only_stripe[5331] = 24'h000000;
assign target_only_stripe[5332] = 24'h000000;
assign target_only_stripe[5333] = 24'h000000;
assign target_only_stripe[5334] = 24'h000000;
assign target_only_stripe[5335] = 24'h000000;
assign target_only_stripe[5336] = 24'h000000;
assign target_only_stripe[5337] = 24'h000000;
assign target_only_stripe[5338] = 24'h000000;
assign target_only_stripe[5339] = 24'h000000;
assign target_only_stripe[5340] = 24'h000000;
assign target_only_stripe[5341] = 24'h000000;
assign target_only_stripe[5342] = 24'h000000;
assign target_only_stripe[5343] = 24'h000000;
assign target_only_stripe[5344] = 24'h000000;
assign target_only_stripe[5345] = 24'h000000;
assign target_only_stripe[5346] = 24'h000000;
assign target_only_stripe[5347] = 24'h000000;
assign target_only_stripe[5348] = 24'h000000;
assign target_only_stripe[5349] = 24'h000000;
assign target_only_stripe[5350] = 24'h000000;
assign target_only_stripe[5351] = 24'h000000;
assign target_only_stripe[5352] = 24'h000000;
assign target_only_stripe[5353] = 24'h000000;
assign target_only_stripe[5354] = 24'h000000;
assign target_only_stripe[5355] = 24'h000000;
assign target_only_stripe[5356] = 24'h000000;
assign target_only_stripe[5357] = 24'h000000;
assign target_only_stripe[5358] = 24'h000000;
assign target_only_stripe[5359] = 24'h000000;
assign target_only_stripe[5360] = 24'h000000;
assign target_only_stripe[5361] = 24'h000000;
assign target_only_stripe[5362] = 24'hffffff;
assign target_only_stripe[5363] = 24'hffffff;
assign target_only_stripe[5364] = 24'hffffff;
assign target_only_stripe[5365] = 24'hffffff;
assign target_only_stripe[5366] = 24'hffffff;
assign target_only_stripe[5367] = 24'hffffff;
assign target_only_stripe[5368] = 24'hffffff;
assign target_only_stripe[5369] = 24'hffffff;
assign target_only_stripe[5370] = 24'hffffff;
assign target_only_stripe[5371] = 24'hffffff;
assign target_only_stripe[5372] = 24'hffffff;
assign target_only_stripe[5373] = 24'hffffff;
assign target_only_stripe[5374] = 24'hffffff;
assign target_only_stripe[5375] = 24'hffffff;
assign target_only_stripe[5376] = 24'hffffff;
assign target_only_stripe[5377] = 24'hffffff;
assign target_only_stripe[5378] = 24'hffffff;
assign target_only_stripe[5379] = 24'hffffff;
assign target_only_stripe[5380] = 24'hffffff;
assign target_only_stripe[5381] = 24'hffffff;
assign target_only_stripe[5382] = 24'hffffff;
assign target_only_stripe[5383] = 24'hffffff;
assign target_only_stripe[5384] = 24'hffffff;
assign target_only_stripe[5385] = 24'hffffff;
assign target_only_stripe[5386] = 24'hffffff;
assign target_only_stripe[5387] = 24'hffffff;
assign target_only_stripe[5388] = 24'hffffff;
assign target_only_stripe[5389] = 24'hffffff;
assign target_only_stripe[5390] = 24'hffffff;
assign target_only_stripe[5391] = 24'hffffff;
assign target_only_stripe[5392] = 24'hffffff;
assign target_only_stripe[5393] = 24'hffffff;
assign target_only_stripe[5394] = 24'hffffff;
assign target_only_stripe[5395] = 24'hffffff;
assign target_only_stripe[5396] = 24'h8e8e8e;
assign target_only_stripe[5397] = 24'h000000;
assign target_only_stripe[5398] = 24'h000000;
assign target_only_stripe[5399] = 24'h000000;
assign target_only_stripe[5400] = 24'h000000;
assign target_only_stripe[5401] = 24'h000000;
assign target_only_stripe[5402] = 24'h000000;
assign target_only_stripe[5403] = 24'h000000;
assign target_only_stripe[5404] = 24'h000000;
assign target_only_stripe[5405] = 24'h000000;
assign target_only_stripe[5406] = 24'h000000;
assign target_only_stripe[5407] = 24'h000000;
assign target_only_stripe[5408] = 24'h000000;
assign target_only_stripe[5409] = 24'h000000;
assign target_only_stripe[5410] = 24'h000000;
assign target_only_stripe[5411] = 24'h000000;
assign target_only_stripe[5412] = 24'h000000;
assign target_only_stripe[5413] = 24'h000000;
assign target_only_stripe[5414] = 24'h000000;
assign target_only_stripe[5415] = 24'h000000;
assign target_only_stripe[5416] = 24'h000000;
assign target_only_stripe[5417] = 24'h000000;
assign target_only_stripe[5418] = 24'h000000;
assign target_only_stripe[5419] = 24'h000000;
assign target_only_stripe[5420] = 24'h000000;
assign target_only_stripe[5421] = 24'h000000;
assign target_only_stripe[5422] = 24'h000000;
assign target_only_stripe[5423] = 24'h000000;
assign target_only_stripe[5424] = 24'h000000;
assign target_only_stripe[5425] = 24'h000000;
assign target_only_stripe[5426] = 24'h000000;
assign target_only_stripe[5427] = 24'h000000;
assign target_only_stripe[5428] = 24'h000000;
assign target_only_stripe[5429] = 24'h000000;
assign target_only_stripe[5430] = 24'h000000;
assign target_only_stripe[5431] = 24'h000000;
assign target_only_stripe[5432] = 24'h000000;
assign target_only_stripe[5433] = 24'h000000;
assign target_only_stripe[5434] = 24'h000000;
assign target_only_stripe[5435] = 24'h000000;
assign target_only_stripe[5436] = 24'h000000;
assign target_only_stripe[5437] = 24'h000000;
assign target_only_stripe[5438] = 24'h000000;
assign target_only_stripe[5439] = 24'h000000;
assign target_only_stripe[5440] = 24'h000000;
assign target_only_stripe[5441] = 24'h000000;
assign target_only_stripe[5442] = 24'h000000;
assign target_only_stripe[5443] = 24'h000000;
assign target_only_stripe[5444] = 24'h000000;
assign target_only_stripe[5445] = 24'h000000;
assign target_only_stripe[5446] = 24'h000000;
assign target_only_stripe[5447] = 24'h000000;
assign target_only_stripe[5448] = 24'h000000;
assign target_only_stripe[5449] = 24'h000000;
assign target_only_stripe[5450] = 24'h000000;
assign target_only_stripe[5451] = 24'h000000;
assign target_only_stripe[5452] = 24'h000000;
assign target_only_stripe[5453] = 24'h000000;
assign target_only_stripe[5454] = 24'h000000;
assign target_only_stripe[5455] = 24'h000000;
assign target_only_stripe[5456] = 24'h000000;
assign target_only_stripe[5457] = 24'h000000;
assign target_only_stripe[5458] = 24'h000000;
assign target_only_stripe[5459] = 24'h000000;
assign target_only_stripe[5460] = 24'hb7b7b7;
assign target_only_stripe[5461] = 24'hffffff;
assign target_only_stripe[5462] = 24'hffffff;
assign target_only_stripe[5463] = 24'hffffff;
assign target_only_stripe[5464] = 24'hffffff;
assign target_only_stripe[5465] = 24'hffffff;
assign target_only_stripe[5466] = 24'hffffff;
assign target_only_stripe[5467] = 24'hffffff;
assign target_only_stripe[5468] = 24'hffffff;
assign target_only_stripe[5469] = 24'hffffff;
assign target_only_stripe[5470] = 24'hffffff;
assign target_only_stripe[5471] = 24'hffffff;
assign target_only_stripe[5472] = 24'hffffff;
assign target_only_stripe[5473] = 24'hffffff;
assign target_only_stripe[5474] = 24'hffffff;
assign target_only_stripe[5475] = 24'hffffff;
assign target_only_stripe[5476] = 24'hffffff;
assign target_only_stripe[5477] = 24'hffffff;
assign target_only_stripe[5478] = 24'hffffff;
assign target_only_stripe[5479] = 24'hffffff;
assign target_only_stripe[5480] = 24'hffffff;
assign target_only_stripe[5481] = 24'hffffff;
assign target_only_stripe[5482] = 24'hffffff;
assign target_only_stripe[5483] = 24'hffffff;
assign target_only_stripe[5484] = 24'hffffff;
assign target_only_stripe[5485] = 24'hffffff;
assign target_only_stripe[5486] = 24'hffffff;
assign target_only_stripe[5487] = 24'hffffff;
assign target_only_stripe[5488] = 24'hffffff;
assign target_only_stripe[5489] = 24'hffffff;
assign target_only_stripe[5490] = 24'hffffff;
assign target_only_stripe[5491] = 24'hffffff;
assign target_only_stripe[5492] = 24'hffffff;
assign target_only_stripe[5493] = 24'hffffff;
assign target_only_stripe[5494] = 24'hefefef;
assign target_only_stripe[5495] = 24'h000000;
assign target_only_stripe[5496] = 24'h000000;
assign target_only_stripe[5497] = 24'h000000;
assign target_only_stripe[5498] = 24'h000000;
assign target_only_stripe[5499] = 24'h000000;
assign target_only_stripe[5500] = 24'h000000;
assign target_only_stripe[5501] = 24'h000000;
assign target_only_stripe[5502] = 24'h000000;
assign target_only_stripe[5503] = 24'h000000;
assign target_only_stripe[5504] = 24'h000000;
assign target_only_stripe[5505] = 24'h000000;
assign target_only_stripe[5506] = 24'h000000;
assign target_only_stripe[5507] = 24'h000000;
assign target_only_stripe[5508] = 24'h000000;
assign target_only_stripe[5509] = 24'h000000;
assign target_only_stripe[5510] = 24'h000000;
assign target_only_stripe[5511] = 24'h000000;
assign target_only_stripe[5512] = 24'h000000;
assign target_only_stripe[5513] = 24'h000000;
assign target_only_stripe[5514] = 24'h000000;
assign target_only_stripe[5515] = 24'h000000;
assign target_only_stripe[5516] = 24'h000000;
assign target_only_stripe[5517] = 24'h000000;
assign target_only_stripe[5518] = 24'h000000;
assign target_only_stripe[5519] = 24'h000000;
assign target_only_stripe[5520] = 24'h000000;
assign target_only_stripe[5521] = 24'h000000;
assign target_only_stripe[5522] = 24'h000000;
assign target_only_stripe[5523] = 24'h000000;
assign target_only_stripe[5524] = 24'h000000;
assign target_only_stripe[5525] = 24'h000000;
assign target_only_stripe[5526] = 24'h000000;
assign target_only_stripe[5527] = 24'hc3c3c3;
assign target_only_stripe[5528] = 24'hffffff;
assign target_only_stripe[5529] = 24'hffffff;
assign target_only_stripe[5530] = 24'hffffff;
assign target_only_stripe[5531] = 24'hffffff;
assign target_only_stripe[5532] = 24'hffffff;
assign target_only_stripe[5533] = 24'hffffff;
assign target_only_stripe[5534] = 24'hffffff;
assign target_only_stripe[5535] = 24'hffffff;
assign target_only_stripe[5536] = 24'hffffff;
assign target_only_stripe[5537] = 24'hffffff;
assign target_only_stripe[5538] = 24'hffffff;
assign target_only_stripe[5539] = 24'hffffff;
assign target_only_stripe[5540] = 24'hffffff;
assign target_only_stripe[5541] = 24'hffffff;
assign target_only_stripe[5542] = 24'hffffff;
assign target_only_stripe[5543] = 24'hffffff;
assign target_only_stripe[5544] = 24'hffffff;
assign target_only_stripe[5545] = 24'hffffff;
assign target_only_stripe[5546] = 24'hffffff;
assign target_only_stripe[5547] = 24'hffffff;
assign target_only_stripe[5548] = 24'hffffff;
assign target_only_stripe[5549] = 24'hffffff;
assign target_only_stripe[5550] = 24'hffffff;
assign target_only_stripe[5551] = 24'hfaf7f5;
assign target_only_stripe[5552] = 24'hebe6db;
assign target_only_stripe[5553] = 24'hffffff;
assign target_only_stripe[5554] = 24'hffffff;
assign target_only_stripe[5555] = 24'hffffff;
assign target_only_stripe[5556] = 24'hffffff;
assign target_only_stripe[5557] = 24'hffffff;
assign target_only_stripe[5558] = 24'hffffff;
assign target_only_stripe[5559] = 24'hffffff;
assign target_only_stripe[5560] = 24'he9e9e9;
assign target_only_stripe[5561] = 24'h191919;
assign target_only_stripe[5562] = 24'h000000;
assign target_only_stripe[5563] = 24'h000000;
assign target_only_stripe[5564] = 24'h000000;
assign target_only_stripe[5565] = 24'h000000;
assign target_only_stripe[5566] = 24'h000000;
assign target_only_stripe[5567] = 24'h000000;
assign target_only_stripe[5568] = 24'h000000;
assign target_only_stripe[5569] = 24'h000000;
assign target_only_stripe[5570] = 24'h000000;
assign target_only_stripe[5571] = 24'h000000;
assign target_only_stripe[5572] = 24'h000000;
assign target_only_stripe[5573] = 24'h000000;
assign target_only_stripe[5574] = 24'h000000;
assign target_only_stripe[5575] = 24'h000000;
assign target_only_stripe[5576] = 24'h000000;
assign target_only_stripe[5577] = 24'h000000;
assign target_only_stripe[5578] = 24'h000000;
assign target_only_stripe[5579] = 24'h000000;
assign target_only_stripe[5580] = 24'h000000;
assign target_only_stripe[5581] = 24'h000000;
assign target_only_stripe[5582] = 24'h000000;
assign target_only_stripe[5583] = 24'h000000;
assign target_only_stripe[5584] = 24'h000000;
assign target_only_stripe[5585] = 24'h000000;
assign target_only_stripe[5586] = 24'h000000;
assign target_only_stripe[5587] = 24'h000000;
assign target_only_stripe[5588] = 24'h000000;
assign target_only_stripe[5589] = 24'h000000;
assign target_only_stripe[5590] = 24'h000000;
assign target_only_stripe[5591] = 24'h000000;
assign target_only_stripe[5592] = 24'h000000;
assign target_only_stripe[5593] = 24'h000000;
assign target_only_stripe[5594] = 24'h000000;
assign target_only_stripe[5595] = 24'h000000;
assign target_only_stripe[5596] = 24'h000000;
assign target_only_stripe[5597] = 24'h000000;
assign target_only_stripe[5598] = 24'h000000;
assign target_only_stripe[5599] = 24'h000000;
assign target_only_stripe[5600] = 24'h000000;
assign target_only_stripe[5601] = 24'h000000;
assign target_only_stripe[5602] = 24'h000000;
assign target_only_stripe[5603] = 24'h000000;
assign target_only_stripe[5604] = 24'h000000;
assign target_only_stripe[5605] = 24'h000000;
assign target_only_stripe[5606] = 24'h000000;
assign target_only_stripe[5607] = 24'h000000;
assign target_only_stripe[5608] = 24'h000000;
assign target_only_stripe[5609] = 24'h000000;
assign target_only_stripe[5610] = 24'h000000;
assign target_only_stripe[5611] = 24'h000000;
assign target_only_stripe[5612] = 24'h000000;
assign target_only_stripe[5613] = 24'h000000;
assign target_only_stripe[5614] = 24'h000000;
assign target_only_stripe[5615] = 24'h000000;
assign target_only_stripe[5616] = 24'h000000;
assign target_only_stripe[5617] = 24'h000000;
assign target_only_stripe[5618] = 24'h000000;
assign target_only_stripe[5619] = 24'h000000;
assign target_only_stripe[5620] = 24'h000000;
assign target_only_stripe[5621] = 24'h000000;
assign target_only_stripe[5622] = 24'h000000;
assign target_only_stripe[5623] = 24'h000000;
assign target_only_stripe[5624] = 24'h0d0d0d;
assign target_only_stripe[5625] = 24'hdcdcdc;
assign target_only_stripe[5626] = 24'hffffff;
assign target_only_stripe[5627] = 24'hffffff;
assign target_only_stripe[5628] = 24'hffffff;
assign target_only_stripe[5629] = 24'hffffff;
assign target_only_stripe[5630] = 24'hffffff;
assign target_only_stripe[5631] = 24'hffffff;
assign target_only_stripe[5632] = 24'hffffff;
assign target_only_stripe[5633] = 24'hffffff;
assign target_only_stripe[5634] = 24'hffffff;
assign target_only_stripe[5635] = 24'hffffff;
assign target_only_stripe[5636] = 24'hffffff;
assign target_only_stripe[5637] = 24'hffffff;
assign target_only_stripe[5638] = 24'hffffff;
assign target_only_stripe[5639] = 24'hffffff;
assign target_only_stripe[5640] = 24'hffffff;
assign target_only_stripe[5641] = 24'hffffff;
assign target_only_stripe[5642] = 24'hffffff;
assign target_only_stripe[5643] = 24'hffffff;
assign target_only_stripe[5644] = 24'hffffff;
assign target_only_stripe[5645] = 24'hffffff;
assign target_only_stripe[5646] = 24'hffffff;
assign target_only_stripe[5647] = 24'hffffff;
assign target_only_stripe[5648] = 24'hffffff;
assign target_only_stripe[5649] = 24'hffffff;
assign target_only_stripe[5650] = 24'hffffff;
assign target_only_stripe[5651] = 24'hffffff;
assign target_only_stripe[5652] = 24'hffffff;
assign target_only_stripe[5653] = 24'hffffff;
assign target_only_stripe[5654] = 24'hffffff;
assign target_only_stripe[5655] = 24'hffffff;
assign target_only_stripe[5656] = 24'hffffff;
assign target_only_stripe[5657] = 24'hffffff;
assign target_only_stripe[5658] = 24'hcccccc;
assign target_only_stripe[5659] = 24'h040404;
assign target_only_stripe[5660] = 24'h000000;
assign target_only_stripe[5661] = 24'h000000;
assign target_only_stripe[5662] = 24'h000000;
assign target_only_stripe[5663] = 24'h000000;
assign target_only_stripe[5664] = 24'h000000;
assign target_only_stripe[5665] = 24'h000000;
assign target_only_stripe[5666] = 24'h000000;
assign target_only_stripe[5667] = 24'h000000;
assign target_only_stripe[5668] = 24'h000000;
assign target_only_stripe[5669] = 24'h000000;
assign target_only_stripe[5670] = 24'h000000;
assign target_only_stripe[5671] = 24'h000000;
assign target_only_stripe[5672] = 24'h000000;
assign target_only_stripe[5673] = 24'h000000;
assign target_only_stripe[5674] = 24'h000000;
assign target_only_stripe[5675] = 24'h000000;
assign target_only_stripe[5676] = 24'h000000;
assign target_only_stripe[5677] = 24'h000000;
assign target_only_stripe[5678] = 24'h000000;
assign target_only_stripe[5679] = 24'h000000;
assign target_only_stripe[5680] = 24'h000000;
assign target_only_stripe[5681] = 24'h000000;
assign target_only_stripe[5682] = 24'h000000;
assign target_only_stripe[5683] = 24'h000000;
assign target_only_stripe[5684] = 24'h000000;
assign target_only_stripe[5685] = 24'h000000;
assign target_only_stripe[5686] = 24'h000000;
assign target_only_stripe[5687] = 24'h000000;
assign target_only_stripe[5688] = 24'h000000;
assign target_only_stripe[5689] = 24'h000000;
assign target_only_stripe[5690] = 24'h000000;
assign target_only_stripe[5691] = 24'hffffff;
assign target_only_stripe[5692] = 24'hffffff;
assign target_only_stripe[5693] = 24'hffffff;
assign target_only_stripe[5694] = 24'hffffff;
assign target_only_stripe[5695] = 24'hffffff;
assign target_only_stripe[5696] = 24'hffffff;
assign target_only_stripe[5697] = 24'hffffff;
assign target_only_stripe[5698] = 24'hffffff;
assign target_only_stripe[5699] = 24'hffffff;
assign target_only_stripe[5700] = 24'hffffff;
assign target_only_stripe[5701] = 24'hffffff;
assign target_only_stripe[5702] = 24'hffffff;
assign target_only_stripe[5703] = 24'hffffff;
assign target_only_stripe[5704] = 24'hffffff;
assign target_only_stripe[5705] = 24'hffffff;
assign target_only_stripe[5706] = 24'hffffff;
assign target_only_stripe[5707] = 24'hffffff;
assign target_only_stripe[5708] = 24'hffffff;
assign target_only_stripe[5709] = 24'hffffff;
assign target_only_stripe[5710] = 24'hffffff;
assign target_only_stripe[5711] = 24'hffffff;
assign target_only_stripe[5712] = 24'hffffff;
assign target_only_stripe[5713] = 24'hffffff;
assign target_only_stripe[5714] = 24'hffffff;
assign target_only_stripe[5715] = 24'hffffff;
assign target_only_stripe[5716] = 24'hffffff;
assign target_only_stripe[5717] = 24'hffffff;
assign target_only_stripe[5718] = 24'hffffff;
assign target_only_stripe[5719] = 24'hffffff;
assign target_only_stripe[5720] = 24'hffffff;
assign target_only_stripe[5721] = 24'hffffff;
assign target_only_stripe[5722] = 24'hffffff;
assign target_only_stripe[5723] = 24'hffffff;
assign target_only_stripe[5724] = 24'hffffff;
assign target_only_stripe[5725] = 24'hadadad;
assign target_only_stripe[5726] = 24'h000000;
assign target_only_stripe[5727] = 24'h000000;
assign target_only_stripe[5728] = 24'h000000;
assign target_only_stripe[5729] = 24'h000000;
assign target_only_stripe[5730] = 24'h000000;
assign target_only_stripe[5731] = 24'h000000;
assign target_only_stripe[5732] = 24'h000000;
assign target_only_stripe[5733] = 24'h000000;
assign target_only_stripe[5734] = 24'h000000;
assign target_only_stripe[5735] = 24'h000000;
assign target_only_stripe[5736] = 24'h000000;
assign target_only_stripe[5737] = 24'h000000;
assign target_only_stripe[5738] = 24'h000000;
assign target_only_stripe[5739] = 24'h000000;
assign target_only_stripe[5740] = 24'h000000;
assign target_only_stripe[5741] = 24'h000000;
assign target_only_stripe[5742] = 24'h000000;
assign target_only_stripe[5743] = 24'h000000;
assign target_only_stripe[5744] = 24'h000000;
assign target_only_stripe[5745] = 24'h000000;
assign target_only_stripe[5746] = 24'h000000;
assign target_only_stripe[5747] = 24'h000000;
assign target_only_stripe[5748] = 24'h000000;
assign target_only_stripe[5749] = 24'h000000;
assign target_only_stripe[5750] = 24'h000000;
assign target_only_stripe[5751] = 24'h000000;
assign target_only_stripe[5752] = 24'h000000;
assign target_only_stripe[5753] = 24'h000000;
assign target_only_stripe[5754] = 24'h000000;
assign target_only_stripe[5755] = 24'h000000;
assign target_only_stripe[5756] = 24'h000000;
assign target_only_stripe[5757] = 24'h000000;
assign target_only_stripe[5758] = 24'h000000;
assign target_only_stripe[5759] = 24'h000000;
assign target_only_stripe[5760] = 24'h000000;
assign target_only_stripe[5761] = 24'h000000;
assign target_only_stripe[5762] = 24'h000000;
assign target_only_stripe[5763] = 24'h000000;
assign target_only_stripe[5764] = 24'h000000;
assign target_only_stripe[5765] = 24'h000000;
assign target_only_stripe[5766] = 24'h000000;
assign target_only_stripe[5767] = 24'h000000;
assign target_only_stripe[5768] = 24'h000000;
assign target_only_stripe[5769] = 24'h000000;
assign target_only_stripe[5770] = 24'h000000;
assign target_only_stripe[5771] = 24'h000000;
assign target_only_stripe[5772] = 24'h000000;
assign target_only_stripe[5773] = 24'h000000;
assign target_only_stripe[5774] = 24'h000000;
assign target_only_stripe[5775] = 24'h000000;
assign target_only_stripe[5776] = 24'h000000;
assign target_only_stripe[5777] = 24'h000000;
assign target_only_stripe[5778] = 24'h000000;
assign target_only_stripe[5779] = 24'h000000;
assign target_only_stripe[5780] = 24'h000000;
assign target_only_stripe[5781] = 24'h000000;
assign target_only_stripe[5782] = 24'h000000;
assign target_only_stripe[5783] = 24'h000000;
assign target_only_stripe[5784] = 24'h000000;
assign target_only_stripe[5785] = 24'h000000;
assign target_only_stripe[5786] = 24'h000000;
assign target_only_stripe[5787] = 24'h000000;
assign target_only_stripe[5788] = 24'h000000;
assign target_only_stripe[5789] = 24'ha7a7a7;
assign target_only_stripe[5790] = 24'hffffff;
assign target_only_stripe[5791] = 24'hffffff;
assign target_only_stripe[5792] = 24'hffffff;
assign target_only_stripe[5793] = 24'hffffff;
assign target_only_stripe[5794] = 24'hffffff;
assign target_only_stripe[5795] = 24'hffffff;
assign target_only_stripe[5796] = 24'hffffff;
assign target_only_stripe[5797] = 24'hffffff;
assign target_only_stripe[5798] = 24'hffffff;
assign target_only_stripe[5799] = 24'hffffff;
assign target_only_stripe[5800] = 24'hffffff;
assign target_only_stripe[5801] = 24'hffffff;
assign target_only_stripe[5802] = 24'hffffff;
assign target_only_stripe[5803] = 24'hffffff;
assign target_only_stripe[5804] = 24'hffffff;
assign target_only_stripe[5805] = 24'hffffff;
assign target_only_stripe[5806] = 24'hffffff;
assign target_only_stripe[5807] = 24'hffffff;
assign target_only_stripe[5808] = 24'hffffff;
assign target_only_stripe[5809] = 24'hffffff;
assign target_only_stripe[5810] = 24'hffffff;
assign target_only_stripe[5811] = 24'hffffff;
assign target_only_stripe[5812] = 24'hffffff;
assign target_only_stripe[5813] = 24'hffffff;
assign target_only_stripe[5814] = 24'hffffff;
assign target_only_stripe[5815] = 24'hffffff;
assign target_only_stripe[5816] = 24'hffffff;
assign target_only_stripe[5817] = 24'hffffff;
assign target_only_stripe[5818] = 24'hffffff;
assign target_only_stripe[5819] = 24'hffffff;
assign target_only_stripe[5820] = 24'hffffff;
assign target_only_stripe[5821] = 24'hffffff;
assign target_only_stripe[5822] = 24'hffffff;
assign target_only_stripe[5823] = 24'hffffff;
assign target_only_stripe[5824] = 24'h000000;
assign target_only_stripe[5825] = 24'h000000;
assign target_only_stripe[5826] = 24'h000000;
assign target_only_stripe[5827] = 24'h000000;
assign target_only_stripe[5828] = 24'h000000;
assign target_only_stripe[5829] = 24'h000000;
assign target_only_stripe[5830] = 24'h000000;
assign target_only_stripe[5831] = 24'h000000;
assign target_only_stripe[5832] = 24'h000000;
assign target_only_stripe[5833] = 24'h000000;
assign target_only_stripe[5834] = 24'h000000;
assign target_only_stripe[5835] = 24'h000000;
assign target_only_stripe[5836] = 24'h000000;
assign target_only_stripe[5837] = 24'h000000;
assign target_only_stripe[5838] = 24'h000000;
assign target_only_stripe[5839] = 24'h000000;
assign target_only_stripe[5840] = 24'h000000;
assign target_only_stripe[5841] = 24'h000000;
assign target_only_stripe[5842] = 24'h000000;
assign target_only_stripe[5843] = 24'h000000;
assign target_only_stripe[5844] = 24'h000000;
assign target_only_stripe[5845] = 24'h000000;
assign target_only_stripe[5846] = 24'h000000;
assign target_only_stripe[5847] = 24'h000000;
assign target_only_stripe[5848] = 24'h000000;
assign target_only_stripe[5849] = 24'h000000;
assign target_only_stripe[5850] = 24'h000000;
assign target_only_stripe[5851] = 24'h000000;
assign target_only_stripe[5852] = 24'h000000;
assign target_only_stripe[5853] = 24'h000000;
assign target_only_stripe[5854] = 24'h000000;
assign target_only_stripe[5855] = 24'h020202;
assign target_only_stripe[5856] = 24'hc7c7c7;
assign target_only_stripe[5857] = 24'hffffff;
assign target_only_stripe[5858] = 24'hffffff;
assign target_only_stripe[5859] = 24'hffffff;
assign target_only_stripe[5860] = 24'hffffff;
assign target_only_stripe[5861] = 24'hffffff;
assign target_only_stripe[5862] = 24'hffffff;
assign target_only_stripe[5863] = 24'hffffff;
assign target_only_stripe[5864] = 24'hffffff;
assign target_only_stripe[5865] = 24'hffffff;
assign target_only_stripe[5866] = 24'hffffff;
assign target_only_stripe[5867] = 24'hffffff;
assign target_only_stripe[5868] = 24'hffffff;
assign target_only_stripe[5869] = 24'hffffff;
assign target_only_stripe[5870] = 24'hffffff;
assign target_only_stripe[5871] = 24'hffffff;
assign target_only_stripe[5872] = 24'hffffff;
assign target_only_stripe[5873] = 24'hffffff;
assign target_only_stripe[5874] = 24'hffffff;
assign target_only_stripe[5875] = 24'hffffff;
assign target_only_stripe[5876] = 24'hffffff;
assign target_only_stripe[5877] = 24'hffffff;
assign target_only_stripe[5878] = 24'hffffff;
assign target_only_stripe[5879] = 24'hffffff;
assign target_only_stripe[5880] = 24'hffffff;
assign target_only_stripe[5881] = 24'hebe6db;
assign target_only_stripe[5882] = 24'hffffff;
assign target_only_stripe[5883] = 24'hfaf7f5;
assign target_only_stripe[5884] = 24'hffffff;
assign target_only_stripe[5885] = 24'hffffff;
assign target_only_stripe[5886] = 24'hffffff;
assign target_only_stripe[5887] = 24'hffffff;
assign target_only_stripe[5888] = 24'hffffff;
assign target_only_stripe[5889] = 24'he1e1e1;
assign target_only_stripe[5890] = 24'h151515;
assign target_only_stripe[5891] = 24'h000000;
assign target_only_stripe[5892] = 24'h000000;
assign target_only_stripe[5893] = 24'h000000;
assign target_only_stripe[5894] = 24'h000000;
assign target_only_stripe[5895] = 24'h000000;
assign target_only_stripe[5896] = 24'h000000;
assign target_only_stripe[5897] = 24'h000000;
assign target_only_stripe[5898] = 24'h000000;
assign target_only_stripe[5899] = 24'h000000;
assign target_only_stripe[5900] = 24'h000000;
assign target_only_stripe[5901] = 24'h000000;
assign target_only_stripe[5902] = 24'h000000;
assign target_only_stripe[5903] = 24'h000000;
assign target_only_stripe[5904] = 24'h000000;
assign target_only_stripe[5905] = 24'h000000;
assign target_only_stripe[5906] = 24'h000000;
assign target_only_stripe[5907] = 24'h000000;
assign target_only_stripe[5908] = 24'h000000;
assign target_only_stripe[5909] = 24'h000000;
assign target_only_stripe[5910] = 24'h000000;
assign target_only_stripe[5911] = 24'h000000;
assign target_only_stripe[5912] = 24'h000000;
assign target_only_stripe[5913] = 24'h000000;
assign target_only_stripe[5914] = 24'h000000;
assign target_only_stripe[5915] = 24'h000000;
assign target_only_stripe[5916] = 24'h000000;
assign target_only_stripe[5917] = 24'h000000;
assign target_only_stripe[5918] = 24'h000000;
assign target_only_stripe[5919] = 24'h000000;
assign target_only_stripe[5920] = 24'h000000;
assign target_only_stripe[5921] = 24'h000000;
assign target_only_stripe[5922] = 24'h000000;
assign target_only_stripe[5923] = 24'h000000;
assign target_only_stripe[5924] = 24'h000000;
assign target_only_stripe[5925] = 24'h000000;
assign target_only_stripe[5926] = 24'h000000;
assign target_only_stripe[5927] = 24'h000000;
assign target_only_stripe[5928] = 24'h000000;
assign target_only_stripe[5929] = 24'h000000;
assign target_only_stripe[5930] = 24'h000000;
assign target_only_stripe[5931] = 24'h000000;
assign target_only_stripe[5932] = 24'h000000;
assign target_only_stripe[5933] = 24'h000000;
assign target_only_stripe[5934] = 24'h000000;
assign target_only_stripe[5935] = 24'h000000;
assign target_only_stripe[5936] = 24'h000000;
assign target_only_stripe[5937] = 24'h000000;
assign target_only_stripe[5938] = 24'h000000;
assign target_only_stripe[5939] = 24'h000000;
assign target_only_stripe[5940] = 24'h000000;
assign target_only_stripe[5941] = 24'h000000;
assign target_only_stripe[5942] = 24'h000000;
assign target_only_stripe[5943] = 24'h000000;
assign target_only_stripe[5944] = 24'h000000;
assign target_only_stripe[5945] = 24'h000000;
assign target_only_stripe[5946] = 24'h000000;
assign target_only_stripe[5947] = 24'h000000;
assign target_only_stripe[5948] = 24'h000000;
assign target_only_stripe[5949] = 24'h000000;
assign target_only_stripe[5950] = 24'h000000;
assign target_only_stripe[5951] = 24'h000000;
assign target_only_stripe[5952] = 24'h000000;
assign target_only_stripe[5953] = 24'h080808;
assign target_only_stripe[5954] = 24'hcfcfcf;
assign target_only_stripe[5955] = 24'hffffff;
assign target_only_stripe[5956] = 24'hffffff;
assign target_only_stripe[5957] = 24'hffffff;
assign target_only_stripe[5958] = 24'hffffff;
assign target_only_stripe[5959] = 24'hffffff;
assign target_only_stripe[5960] = 24'hffffff;
assign target_only_stripe[5961] = 24'hffffff;
assign target_only_stripe[5962] = 24'hffffff;
assign target_only_stripe[5963] = 24'hffffff;
assign target_only_stripe[5964] = 24'hffffff;
assign target_only_stripe[5965] = 24'hffffff;
assign target_only_stripe[5966] = 24'hffffff;
assign target_only_stripe[5967] = 24'hffffff;
assign target_only_stripe[5968] = 24'hffffff;
assign target_only_stripe[5969] = 24'hffffff;
assign target_only_stripe[5970] = 24'hffffff;
assign target_only_stripe[5971] = 24'hffffff;
assign target_only_stripe[5972] = 24'hffffff;
assign target_only_stripe[5973] = 24'hffffff;
assign target_only_stripe[5974] = 24'hffffff;
assign target_only_stripe[5975] = 24'hffffff;
assign target_only_stripe[5976] = 24'hffffff;
assign target_only_stripe[5977] = 24'hffffff;
assign target_only_stripe[5978] = 24'hffffff;
assign target_only_stripe[5979] = 24'hffffff;
assign target_only_stripe[5980] = 24'hffffff;
assign target_only_stripe[5981] = 24'hffffff;
assign target_only_stripe[5982] = 24'hffffff;
assign target_only_stripe[5983] = 24'hffffff;
assign target_only_stripe[5984] = 24'hffffff;
assign target_only_stripe[5985] = 24'hffffff;
assign target_only_stripe[5986] = 24'hffffff;
assign target_only_stripe[5987] = 24'hd2d2d2;
assign target_only_stripe[5988] = 24'h0e0e0e;
assign target_only_stripe[5989] = 24'h000000;
assign target_only_stripe[5990] = 24'h000000;
assign target_only_stripe[5991] = 24'h000000;
assign target_only_stripe[5992] = 24'h000000;
assign target_only_stripe[5993] = 24'h000000;
assign target_only_stripe[5994] = 24'h000000;
assign target_only_stripe[5995] = 24'h000000;
assign target_only_stripe[5996] = 24'h000000;
assign target_only_stripe[5997] = 24'h000000;
assign target_only_stripe[5998] = 24'h000000;
assign target_only_stripe[5999] = 24'h000000;
assign target_only_stripe[6000] = 24'h000000;
assign target_only_stripe[6001] = 24'h000000;
assign target_only_stripe[6002] = 24'h000000;
assign target_only_stripe[6003] = 24'h000000;
assign target_only_stripe[6004] = 24'h000000;
assign target_only_stripe[6005] = 24'h000000;
assign target_only_stripe[6006] = 24'h000000;
assign target_only_stripe[6007] = 24'h000000;
assign target_only_stripe[6008] = 24'h000000;
assign target_only_stripe[6009] = 24'h000000;
assign target_only_stripe[6010] = 24'h000000;
assign target_only_stripe[6011] = 24'h000000;
assign target_only_stripe[6012] = 24'h000000;
assign target_only_stripe[6013] = 24'h000000;
assign target_only_stripe[6014] = 24'h000000;
assign target_only_stripe[6015] = 24'h000000;
assign target_only_stripe[6016] = 24'h000000;
assign target_only_stripe[6017] = 24'h000000;
assign target_only_stripe[6018] = 24'h000000;
assign target_only_stripe[6019] = 24'h000000;
assign target_only_stripe[6020] = 24'h3a3a3a;
assign target_only_stripe[6021] = 24'hffffff;
assign target_only_stripe[6022] = 24'hffffff;
assign target_only_stripe[6023] = 24'hffffff;
assign target_only_stripe[6024] = 24'hffffff;
assign target_only_stripe[6025] = 24'hffffff;
assign target_only_stripe[6026] = 24'hffffff;
assign target_only_stripe[6027] = 24'hffffff;
assign target_only_stripe[6028] = 24'hffffff;
assign target_only_stripe[6029] = 24'hffffff;
assign target_only_stripe[6030] = 24'hffffff;
assign target_only_stripe[6031] = 24'hffffff;
assign target_only_stripe[6032] = 24'hffffff;
assign target_only_stripe[6033] = 24'hffffff;
assign target_only_stripe[6034] = 24'hffffff;
assign target_only_stripe[6035] = 24'hffffff;
assign target_only_stripe[6036] = 24'hffffff;
assign target_only_stripe[6037] = 24'hffffff;
assign target_only_stripe[6038] = 24'hffffff;
assign target_only_stripe[6039] = 24'hffffff;
assign target_only_stripe[6040] = 24'hffffff;
assign target_only_stripe[6041] = 24'hffffff;
assign target_only_stripe[6042] = 24'hffffff;
assign target_only_stripe[6043] = 24'hffffff;
assign target_only_stripe[6044] = 24'hffffff;
assign target_only_stripe[6045] = 24'hffffff;
assign target_only_stripe[6046] = 24'hffffff;
assign target_only_stripe[6047] = 24'hffffff;
assign target_only_stripe[6048] = 24'hffffff;
assign target_only_stripe[6049] = 24'hffffff;
assign target_only_stripe[6050] = 24'hffffff;
assign target_only_stripe[6051] = 24'hffffff;
assign target_only_stripe[6052] = 24'hffffff;
assign target_only_stripe[6053] = 24'hffffff;
assign target_only_stripe[6054] = 24'hffffff;
assign target_only_stripe[6055] = 24'h0b0b0b;
assign target_only_stripe[6056] = 24'h000000;
assign target_only_stripe[6057] = 24'h000000;
assign target_only_stripe[6058] = 24'h000000;
assign target_only_stripe[6059] = 24'h000000;
assign target_only_stripe[6060] = 24'h000000;
assign target_only_stripe[6061] = 24'h000000;
assign target_only_stripe[6062] = 24'h000000;
assign target_only_stripe[6063] = 24'h000000;
assign target_only_stripe[6064] = 24'h000000;
assign target_only_stripe[6065] = 24'h000000;
assign target_only_stripe[6066] = 24'h000000;
assign target_only_stripe[6067] = 24'h000000;
assign target_only_stripe[6068] = 24'h000000;
assign target_only_stripe[6069] = 24'h000000;
assign target_only_stripe[6070] = 24'h000000;
assign target_only_stripe[6071] = 24'h000000;
assign target_only_stripe[6072] = 24'h000000;
assign target_only_stripe[6073] = 24'h000000;
assign target_only_stripe[6074] = 24'h000000;
assign target_only_stripe[6075] = 24'h000000;
assign target_only_stripe[6076] = 24'h000000;
assign target_only_stripe[6077] = 24'h000000;
assign target_only_stripe[6078] = 24'h000000;
assign target_only_stripe[6079] = 24'h000000;
assign target_only_stripe[6080] = 24'h000000;
assign target_only_stripe[6081] = 24'h000000;
assign target_only_stripe[6082] = 24'h000000;
assign target_only_stripe[6083] = 24'h000000;
assign target_only_stripe[6084] = 24'h000000;
assign target_only_stripe[6085] = 24'h000000;
assign target_only_stripe[6086] = 24'h000000;
assign target_only_stripe[6087] = 24'h000000;
assign target_only_stripe[6088] = 24'h000000;
assign target_only_stripe[6089] = 24'h000000;
assign target_only_stripe[6090] = 24'h000000;
assign target_only_stripe[6091] = 24'h000000;
assign target_only_stripe[6092] = 24'h000000;
assign target_only_stripe[6093] = 24'h000000;
assign target_only_stripe[6094] = 24'h000000;
assign target_only_stripe[6095] = 24'h000000;
assign target_only_stripe[6096] = 24'h000000;
assign target_only_stripe[6097] = 24'h000000;
assign target_only_stripe[6098] = 24'h000000;
assign target_only_stripe[6099] = 24'h000000;
assign target_only_stripe[6100] = 24'h000000;
assign target_only_stripe[6101] = 24'h000000;
assign target_only_stripe[6102] = 24'h000000;
assign target_only_stripe[6103] = 24'h000000;
assign target_only_stripe[6104] = 24'h000000;
assign target_only_stripe[6105] = 24'h000000;
assign target_only_stripe[6106] = 24'h000000;
assign target_only_stripe[6107] = 24'h000000;
assign target_only_stripe[6108] = 24'h000000;
assign target_only_stripe[6109] = 24'h000000;
assign target_only_stripe[6110] = 24'h000000;
assign target_only_stripe[6111] = 24'h000000;
assign target_only_stripe[6112] = 24'h000000;
assign target_only_stripe[6113] = 24'h000000;
assign target_only_stripe[6114] = 24'h000000;
assign target_only_stripe[6115] = 24'h000000;
assign target_only_stripe[6116] = 24'h000000;
assign target_only_stripe[6117] = 24'h080808;
assign target_only_stripe[6118] = 24'hffffff;
assign target_only_stripe[6119] = 24'hffffff;
assign target_only_stripe[6120] = 24'hffffff;
assign target_only_stripe[6121] = 24'hffffff;
assign target_only_stripe[6122] = 24'hffffff;
assign target_only_stripe[6123] = 24'hffffff;
assign target_only_stripe[6124] = 24'hffffff;
assign target_only_stripe[6125] = 24'hffffff;
assign target_only_stripe[6126] = 24'hffffff;
assign target_only_stripe[6127] = 24'hffffff;
assign target_only_stripe[6128] = 24'hffffff;
assign target_only_stripe[6129] = 24'hffffff;
assign target_only_stripe[6130] = 24'hffffff;
assign target_only_stripe[6131] = 24'hffffff;
assign target_only_stripe[6132] = 24'hffffff;
assign target_only_stripe[6133] = 24'hffffff;
assign target_only_stripe[6134] = 24'hffffff;
assign target_only_stripe[6135] = 24'hffffff;
assign target_only_stripe[6136] = 24'hffffff;
assign target_only_stripe[6137] = 24'hffffff;
assign target_only_stripe[6138] = 24'hffffff;
assign target_only_stripe[6139] = 24'hffffff;
assign target_only_stripe[6140] = 24'hffffff;
assign target_only_stripe[6141] = 24'hffffff;
assign target_only_stripe[6142] = 24'hffffff;
assign target_only_stripe[6143] = 24'hffffff;
assign target_only_stripe[6144] = 24'hffffff;
assign target_only_stripe[6145] = 24'hffffff;
assign target_only_stripe[6146] = 24'hffffff;
assign target_only_stripe[6147] = 24'hffffff;
assign target_only_stripe[6148] = 24'hffffff;
assign target_only_stripe[6149] = 24'hffffff;
assign target_only_stripe[6150] = 24'hffffff;
assign target_only_stripe[6151] = 24'hffffff;
assign target_only_stripe[6152] = 24'h454545;
assign target_only_stripe[6153] = 24'h000000;
assign target_only_stripe[6154] = 24'h000000;
assign target_only_stripe[6155] = 24'h000000;
assign target_only_stripe[6156] = 24'h000000;
assign target_only_stripe[6157] = 24'h000000;
assign target_only_stripe[6158] = 24'h000000;
assign target_only_stripe[6159] = 24'h000000;
assign target_only_stripe[6160] = 24'h000000;
assign target_only_stripe[6161] = 24'h000000;
assign target_only_stripe[6162] = 24'h000000;
assign target_only_stripe[6163] = 24'h000000;
assign target_only_stripe[6164] = 24'h000000;
assign target_only_stripe[6165] = 24'h000000;
assign target_only_stripe[6166] = 24'h000000;
assign target_only_stripe[6167] = 24'h000000;
assign target_only_stripe[6168] = 24'h000000;
assign target_only_stripe[6169] = 24'h000000;
assign target_only_stripe[6170] = 24'h000000;
assign target_only_stripe[6171] = 24'h000000;
assign target_only_stripe[6172] = 24'h000000;
assign target_only_stripe[6173] = 24'h000000;
assign target_only_stripe[6174] = 24'h000000;
assign target_only_stripe[6175] = 24'h000000;
assign target_only_stripe[6176] = 24'h000000;
assign target_only_stripe[6177] = 24'h000000;
assign target_only_stripe[6178] = 24'h000000;
assign target_only_stripe[6179] = 24'h000000;
assign target_only_stripe[6180] = 24'h000000;
assign target_only_stripe[6181] = 24'h000000;
assign target_only_stripe[6182] = 24'h000000;
assign target_only_stripe[6183] = 24'h000000;
assign target_only_stripe[6184] = 24'h090909;
assign target_only_stripe[6185] = 24'hcdcdcd;
assign target_only_stripe[6186] = 24'hffffff;
assign target_only_stripe[6187] = 24'hffffff;
assign target_only_stripe[6188] = 24'hffffff;
assign target_only_stripe[6189] = 24'hffffff;
assign target_only_stripe[6190] = 24'hffffff;
assign target_only_stripe[6191] = 24'hffffff;
assign target_only_stripe[6192] = 24'hffffff;
assign target_only_stripe[6193] = 24'hffffff;
assign target_only_stripe[6194] = 24'hffffff;
assign target_only_stripe[6195] = 24'hffffff;
assign target_only_stripe[6196] = 24'hffffff;
assign target_only_stripe[6197] = 24'hffffff;
assign target_only_stripe[6198] = 24'hffffff;
assign target_only_stripe[6199] = 24'hffffff;
assign target_only_stripe[6200] = 24'hffffff;
assign target_only_stripe[6201] = 24'hffffff;
assign target_only_stripe[6202] = 24'hffffff;
assign target_only_stripe[6203] = 24'hffffff;
assign target_only_stripe[6204] = 24'hffffff;
assign target_only_stripe[6205] = 24'hffffff;
assign target_only_stripe[6206] = 24'hffffff;
assign target_only_stripe[6207] = 24'hffffff;
assign target_only_stripe[6208] = 24'hffffff;
assign target_only_stripe[6209] = 24'hffffff;
assign target_only_stripe[6210] = 24'hffffff;
assign target_only_stripe[6211] = 24'hffffff;
assign target_only_stripe[6212] = 24'hfaf7f5;
assign target_only_stripe[6213] = 24'hffffff;
assign target_only_stripe[6214] = 24'hffffff;
assign target_only_stripe[6215] = 24'hffffff;
assign target_only_stripe[6216] = 24'hffffff;
assign target_only_stripe[6217] = 24'hffffff;
assign target_only_stripe[6218] = 24'hd4d4d4;
assign target_only_stripe[6219] = 24'h0e0e0e;
assign target_only_stripe[6220] = 24'h000000;
assign target_only_stripe[6221] = 24'h000000;
assign target_only_stripe[6222] = 24'h000000;
assign target_only_stripe[6223] = 24'h000000;
assign target_only_stripe[6224] = 24'h000000;
assign target_only_stripe[6225] = 24'h000000;
assign target_only_stripe[6226] = 24'h000000;
assign target_only_stripe[6227] = 24'h000000;
assign target_only_stripe[6228] = 24'h000000;
assign target_only_stripe[6229] = 24'h000000;
assign target_only_stripe[6230] = 24'h000000;
assign target_only_stripe[6231] = 24'h000000;
assign target_only_stripe[6232] = 24'h000000;
assign target_only_stripe[6233] = 24'h000000;
assign target_only_stripe[6234] = 24'h000000;
assign target_only_stripe[6235] = 24'h000000;
assign target_only_stripe[6236] = 24'h000000;
assign target_only_stripe[6237] = 24'h000000;
assign target_only_stripe[6238] = 24'h000000;
assign target_only_stripe[6239] = 24'h000000;
assign target_only_stripe[6240] = 24'h000000;
assign target_only_stripe[6241] = 24'h000000;
assign target_only_stripe[6242] = 24'h000000;
assign target_only_stripe[6243] = 24'h000000;
assign target_only_stripe[6244] = 24'h000000;
assign target_only_stripe[6245] = 24'h000000;
assign target_only_stripe[6246] = 24'h000000;
assign target_only_stripe[6247] = 24'h000000;
assign target_only_stripe[6248] = 24'h000000;
assign target_only_stripe[6249] = 24'h000000;
assign target_only_stripe[6250] = 24'h000000;
assign target_only_stripe[6251] = 24'h000000;
assign target_only_stripe[6252] = 24'h000000;
assign target_only_stripe[6253] = 24'h000000;
assign target_only_stripe[6254] = 24'h000000;
assign target_only_stripe[6255] = 24'h000000;
assign target_only_stripe[6256] = 24'h000000;
assign target_only_stripe[6257] = 24'h000000;
assign target_only_stripe[6258] = 24'h000000;
assign target_only_stripe[6259] = 24'h000000;
assign target_only_stripe[6260] = 24'h000000;
assign target_only_stripe[6261] = 24'h000000;
assign target_only_stripe[6262] = 24'h000000;
assign target_only_stripe[6263] = 24'h000000;
assign target_only_stripe[6264] = 24'h000000;
assign target_only_stripe[6265] = 24'h000000;
assign target_only_stripe[6266] = 24'h000000;
assign target_only_stripe[6267] = 24'h000000;
assign target_only_stripe[6268] = 24'h000000;
assign target_only_stripe[6269] = 24'h000000;
assign target_only_stripe[6270] = 24'h000000;
assign target_only_stripe[6271] = 24'h000000;
assign target_only_stripe[6272] = 24'h000000;
assign target_only_stripe[6273] = 24'h000000;
assign target_only_stripe[6274] = 24'h000000;
assign target_only_stripe[6275] = 24'h000000;
assign target_only_stripe[6276] = 24'h000000;
assign target_only_stripe[6277] = 24'h000000;
assign target_only_stripe[6278] = 24'h000000;
assign target_only_stripe[6279] = 24'h000000;
assign target_only_stripe[6280] = 24'h000000;
assign target_only_stripe[6281] = 24'h000000;
assign target_only_stripe[6282] = 24'h010101;
assign target_only_stripe[6283] = 24'hbfbfbf;
assign target_only_stripe[6284] = 24'hffffff;
assign target_only_stripe[6285] = 24'hffffff;
assign target_only_stripe[6286] = 24'hffffff;
assign target_only_stripe[6287] = 24'hffffff;
assign target_only_stripe[6288] = 24'hffffff;
assign target_only_stripe[6289] = 24'hffffff;
assign target_only_stripe[6290] = 24'hfaf7f5;
assign target_only_stripe[6291] = 24'hffffff;
assign target_only_stripe[6292] = 24'hffffff;
assign target_only_stripe[6293] = 24'hffffff;
assign target_only_stripe[6294] = 24'hffffff;
assign target_only_stripe[6295] = 24'hffffff;
assign target_only_stripe[6296] = 24'hffffff;
assign target_only_stripe[6297] = 24'hffffff;
assign target_only_stripe[6298] = 24'hffffff;
assign target_only_stripe[6299] = 24'hffffff;
assign target_only_stripe[6300] = 24'hffffff;
assign target_only_stripe[6301] = 24'hffffff;
assign target_only_stripe[6302] = 24'hffffff;
assign target_only_stripe[6303] = 24'hffffff;
assign target_only_stripe[6304] = 24'hffffff;
assign target_only_stripe[6305] = 24'hffffff;
assign target_only_stripe[6306] = 24'hffffff;
assign target_only_stripe[6307] = 24'hffffff;
assign target_only_stripe[6308] = 24'hffffff;
assign target_only_stripe[6309] = 24'hffffff;
assign target_only_stripe[6310] = 24'hffffff;
assign target_only_stripe[6311] = 24'hffffff;
assign target_only_stripe[6312] = 24'hffffff;
assign target_only_stripe[6313] = 24'hffffff;
assign target_only_stripe[6314] = 24'hffffff;
assign target_only_stripe[6315] = 24'hffffff;
assign target_only_stripe[6316] = 24'hdcdcdc;
assign target_only_stripe[6317] = 24'h191919;
assign target_only_stripe[6318] = 24'h000000;
assign target_only_stripe[6319] = 24'h000000;
assign target_only_stripe[6320] = 24'h000000;
assign target_only_stripe[6321] = 24'h000000;
assign target_only_stripe[6322] = 24'h000000;
assign target_only_stripe[6323] = 24'h000000;
assign target_only_stripe[6324] = 24'h000000;
assign target_only_stripe[6325] = 24'h000000;
assign target_only_stripe[6326] = 24'h000000;
assign target_only_stripe[6327] = 24'h000000;
assign target_only_stripe[6328] = 24'h000000;
assign target_only_stripe[6329] = 24'h000000;
assign target_only_stripe[6330] = 24'h000000;
assign target_only_stripe[6331] = 24'h000000;
assign target_only_stripe[6332] = 24'h000000;
assign target_only_stripe[6333] = 24'h000000;
assign target_only_stripe[6334] = 24'h000000;
assign target_only_stripe[6335] = 24'h000000;
assign target_only_stripe[6336] = 24'h000000;
assign target_only_stripe[6337] = 24'h000000;
assign target_only_stripe[6338] = 24'h000000;
assign target_only_stripe[6339] = 24'h000000;
assign target_only_stripe[6340] = 24'h000000;
assign target_only_stripe[6341] = 24'h000000;
assign target_only_stripe[6342] = 24'h000000;
assign target_only_stripe[6343] = 24'h000000;
assign target_only_stripe[6344] = 24'h000000;
assign target_only_stripe[6345] = 24'h000000;
assign target_only_stripe[6346] = 24'h000000;
assign target_only_stripe[6347] = 24'h000000;
assign target_only_stripe[6348] = 24'h000000;
assign target_only_stripe[6349] = 24'h313131;
assign target_only_stripe[6350] = 24'hffffff;
assign target_only_stripe[6351] = 24'hffffff;
assign target_only_stripe[6352] = 24'hffffff;
assign target_only_stripe[6353] = 24'hffffff;
assign target_only_stripe[6354] = 24'hffffff;
assign target_only_stripe[6355] = 24'hffffff;
assign target_only_stripe[6356] = 24'hffffff;
assign target_only_stripe[6357] = 24'hffffff;
assign target_only_stripe[6358] = 24'hffffff;
assign target_only_stripe[6359] = 24'hffffff;
assign target_only_stripe[6360] = 24'hffffff;
assign target_only_stripe[6361] = 24'hffffff;
assign target_only_stripe[6362] = 24'hffffff;
assign target_only_stripe[6363] = 24'hffffff;
assign target_only_stripe[6364] = 24'hffffff;
assign target_only_stripe[6365] = 24'hffffff;
assign target_only_stripe[6366] = 24'hffffff;
assign target_only_stripe[6367] = 24'hffffff;
assign target_only_stripe[6368] = 24'hffffff;
assign target_only_stripe[6369] = 24'hffffff;
assign target_only_stripe[6370] = 24'hffffff;
assign target_only_stripe[6371] = 24'hffffff;
assign target_only_stripe[6372] = 24'hffffff;
assign target_only_stripe[6373] = 24'hffffff;
assign target_only_stripe[6374] = 24'hffffff;
assign target_only_stripe[6375] = 24'hffffff;
assign target_only_stripe[6376] = 24'hffffff;
assign target_only_stripe[6377] = 24'hffffff;
assign target_only_stripe[6378] = 24'hffffff;
assign target_only_stripe[6379] = 24'hffffff;
assign target_only_stripe[6380] = 24'hffffff;
assign target_only_stripe[6381] = 24'hffffff;
assign target_only_stripe[6382] = 24'hffffff;
assign target_only_stripe[6383] = 24'hffffff;
assign target_only_stripe[6384] = 24'h525252;
assign target_only_stripe[6385] = 24'h000000;
assign target_only_stripe[6386] = 24'h000000;
assign target_only_stripe[6387] = 24'h000000;
assign target_only_stripe[6388] = 24'h000000;
assign target_only_stripe[6389] = 24'h000000;
assign target_only_stripe[6390] = 24'h000000;
assign target_only_stripe[6391] = 24'h000000;
assign target_only_stripe[6392] = 24'h000000;
assign target_only_stripe[6393] = 24'h000000;
assign target_only_stripe[6394] = 24'h000000;
assign target_only_stripe[6395] = 24'h000000;
assign target_only_stripe[6396] = 24'h000000;
assign target_only_stripe[6397] = 24'h000000;
assign target_only_stripe[6398] = 24'h000000;
assign target_only_stripe[6399] = 24'h000000;
assign target_only_stripe[6400] = 24'h000000;
assign target_only_stripe[6401] = 24'h000000;
assign target_only_stripe[6402] = 24'h000000;
assign target_only_stripe[6403] = 24'h000000;
assign target_only_stripe[6404] = 24'h000000;
assign target_only_stripe[6405] = 24'h000000;
assign target_only_stripe[6406] = 24'h000000;
assign target_only_stripe[6407] = 24'h000000;
assign target_only_stripe[6408] = 24'h000000;
assign target_only_stripe[6409] = 24'h000000;
assign target_only_stripe[6410] = 24'h000000;
assign target_only_stripe[6411] = 24'h000000;
assign target_only_stripe[6412] = 24'h000000;
assign target_only_stripe[6413] = 24'h000000;
assign target_only_stripe[6414] = 24'h000000;
assign target_only_stripe[6415] = 24'h000000;
assign target_only_stripe[6416] = 24'h000000;
assign target_only_stripe[6417] = 24'h000000;
assign target_only_stripe[6418] = 24'h000000;
assign target_only_stripe[6419] = 24'h000000;
assign target_only_stripe[6420] = 24'h000000;
assign target_only_stripe[6421] = 24'h000000;
assign target_only_stripe[6422] = 24'h000000;
assign target_only_stripe[6423] = 24'h000000;
assign target_only_stripe[6424] = 24'h000000;
assign target_only_stripe[6425] = 24'h000000;
assign target_only_stripe[6426] = 24'h000000;
assign target_only_stripe[6427] = 24'h000000;
assign target_only_stripe[6428] = 24'h000000;
assign target_only_stripe[6429] = 24'h000000;
assign target_only_stripe[6430] = 24'h000000;
assign target_only_stripe[6431] = 24'h000000;
assign target_only_stripe[6432] = 24'h000000;
assign target_only_stripe[6433] = 24'h000000;
assign target_only_stripe[6434] = 24'h000000;
assign target_only_stripe[6435] = 24'h000000;
assign target_only_stripe[6436] = 24'h000000;
assign target_only_stripe[6437] = 24'h000000;
assign target_only_stripe[6438] = 24'h000000;
assign target_only_stripe[6439] = 24'h000000;
assign target_only_stripe[6440] = 24'h000000;
assign target_only_stripe[6441] = 24'h000000;
assign target_only_stripe[6442] = 24'h000000;
assign target_only_stripe[6443] = 24'h000000;
assign target_only_stripe[6444] = 24'h000000;
assign target_only_stripe[6445] = 24'h000000;
assign target_only_stripe[6446] = 24'h424242;
assign target_only_stripe[6447] = 24'hd2c7c4;
assign target_only_stripe[6448] = 24'hffffff;
assign target_only_stripe[6449] = 24'hffffff;
assign target_only_stripe[6450] = 24'hffffff;
assign target_only_stripe[6451] = 24'hffffff;
assign target_only_stripe[6452] = 24'hffffff;
assign target_only_stripe[6453] = 24'hffffff;
assign target_only_stripe[6454] = 24'hffffff;
assign target_only_stripe[6455] = 24'hffffff;
assign target_only_stripe[6456] = 24'hffffff;
assign target_only_stripe[6457] = 24'hffffff;
assign target_only_stripe[6458] = 24'hffffff;
assign target_only_stripe[6459] = 24'hffffff;
assign target_only_stripe[6460] = 24'hffffff;
assign target_only_stripe[6461] = 24'hffffff;
assign target_only_stripe[6462] = 24'hffffff;
assign target_only_stripe[6463] = 24'hffffff;
assign target_only_stripe[6464] = 24'hffffff;
assign target_only_stripe[6465] = 24'hffffff;
assign target_only_stripe[6466] = 24'hffffff;
assign target_only_stripe[6467] = 24'hffffff;
assign target_only_stripe[6468] = 24'hffffff;
assign target_only_stripe[6469] = 24'hffffff;
assign target_only_stripe[6470] = 24'hffffff;
assign target_only_stripe[6471] = 24'hffffff;
assign target_only_stripe[6472] = 24'hffffff;
assign target_only_stripe[6473] = 24'hffffff;
assign target_only_stripe[6474] = 24'hffffff;
assign target_only_stripe[6475] = 24'hffffff;
assign target_only_stripe[6476] = 24'hffffff;
assign target_only_stripe[6477] = 24'hffffff;
assign target_only_stripe[6478] = 24'hffffff;
assign target_only_stripe[6479] = 24'hffffff;
assign target_only_stripe[6480] = 24'hbfb1ab;
assign target_only_stripe[6481] = 24'h3a3a3a;
assign target_only_stripe[6482] = 24'h000000;
assign target_only_stripe[6483] = 24'h000000;
assign target_only_stripe[6484] = 24'h000000;
assign target_only_stripe[6485] = 24'h000000;
assign target_only_stripe[6486] = 24'h000000;
assign target_only_stripe[6487] = 24'h000000;
assign target_only_stripe[6488] = 24'h000000;
assign target_only_stripe[6489] = 24'h000000;
assign target_only_stripe[6490] = 24'h000000;
assign target_only_stripe[6491] = 24'h000000;
assign target_only_stripe[6492] = 24'h000000;
assign target_only_stripe[6493] = 24'h000000;
assign target_only_stripe[6494] = 24'h000000;
assign target_only_stripe[6495] = 24'h000000;
assign target_only_stripe[6496] = 24'h000000;
assign target_only_stripe[6497] = 24'h000000;
assign target_only_stripe[6498] = 24'h000000;
assign target_only_stripe[6499] = 24'h000000;
assign target_only_stripe[6500] = 24'h000000;
assign target_only_stripe[6501] = 24'h000000;
assign target_only_stripe[6502] = 24'h000000;
assign target_only_stripe[6503] = 24'h000000;
assign target_only_stripe[6504] = 24'h000000;
assign target_only_stripe[6505] = 24'h000000;
assign target_only_stripe[6506] = 24'h000000;
assign target_only_stripe[6507] = 24'h000000;
assign target_only_stripe[6508] = 24'h000000;
assign target_only_stripe[6509] = 24'h000000;
assign target_only_stripe[6510] = 24'h000000;
assign target_only_stripe[6511] = 24'h000000;
assign target_only_stripe[6512] = 24'h000000;
assign target_only_stripe[6513] = 24'h121212;
assign target_only_stripe[6514] = 24'hd7d7d7;
assign target_only_stripe[6515] = 24'hffffff;
assign target_only_stripe[6516] = 24'hffffff;
assign target_only_stripe[6517] = 24'hffffff;
assign target_only_stripe[6518] = 24'hffffff;
assign target_only_stripe[6519] = 24'hffffff;
assign target_only_stripe[6520] = 24'hffffff;
assign target_only_stripe[6521] = 24'hffffff;
assign target_only_stripe[6522] = 24'hffffff;
assign target_only_stripe[6523] = 24'hffffff;
assign target_only_stripe[6524] = 24'hffffff;
assign target_only_stripe[6525] = 24'hffffff;
assign target_only_stripe[6526] = 24'hffffff;
assign target_only_stripe[6527] = 24'hffffff;
assign target_only_stripe[6528] = 24'hffffff;
assign target_only_stripe[6529] = 24'hffffff;
assign target_only_stripe[6530] = 24'hffffff;
assign target_only_stripe[6531] = 24'hffffff;
assign target_only_stripe[6532] = 24'hffffff;
assign target_only_stripe[6533] = 24'hffffff;
assign target_only_stripe[6534] = 24'hffffff;
assign target_only_stripe[6535] = 24'hffffff;
assign target_only_stripe[6536] = 24'hffffff;
assign target_only_stripe[6537] = 24'hffffff;
assign target_only_stripe[6538] = 24'hffffff;
assign target_only_stripe[6539] = 24'hffffff;
assign target_only_stripe[6540] = 24'hffffff;
assign target_only_stripe[6541] = 24'hfaf7f5;
assign target_only_stripe[6542] = 24'hffffff;
assign target_only_stripe[6543] = 24'hffffff;
assign target_only_stripe[6544] = 24'hffffff;
assign target_only_stripe[6545] = 24'hffffff;
assign target_only_stripe[6546] = 24'hffffff;
assign target_only_stripe[6547] = 24'hc5c5c5;
assign target_only_stripe[6548] = 24'h030303;
assign target_only_stripe[6549] = 24'h000000;
assign target_only_stripe[6550] = 24'h000000;
assign target_only_stripe[6551] = 24'h000000;
assign target_only_stripe[6552] = 24'h000000;
assign target_only_stripe[6553] = 24'h000000;
assign target_only_stripe[6554] = 24'h000000;
assign target_only_stripe[6555] = 24'h000000;
assign target_only_stripe[6556] = 24'h000000;
assign target_only_stripe[6557] = 24'h000000;
assign target_only_stripe[6558] = 24'h000000;
assign target_only_stripe[6559] = 24'h000000;
assign target_only_stripe[6560] = 24'h000000;
assign target_only_stripe[6561] = 24'h000000;
assign target_only_stripe[6562] = 24'h000000;
assign target_only_stripe[6563] = 24'h000000;
assign target_only_stripe[6564] = 24'h000000;
assign target_only_stripe[6565] = 24'h000000;
assign target_only_stripe[6566] = 24'h000000;
assign target_only_stripe[6567] = 24'h000000;
assign target_only_stripe[6568] = 24'h000000;
assign target_only_stripe[6569] = 24'h000000;
assign target_only_stripe[6570] = 24'h000000;
assign target_only_stripe[6571] = 24'h000000;
assign target_only_stripe[6572] = 24'h000000;
assign target_only_stripe[6573] = 24'h000000;
assign target_only_stripe[6574] = 24'h000000;
assign target_only_stripe[6575] = 24'h000000;
assign target_only_stripe[6576] = 24'h000000;
assign target_only_stripe[6577] = 24'h000000;
assign target_only_stripe[6578] = 24'h000000;
assign target_only_stripe[6579] = 24'h000000;
assign target_only_stripe[6580] = 24'h000000;
assign target_only_stripe[6581] = 24'h000000;
assign target_only_stripe[6582] = 24'h000000;
assign target_only_stripe[6583] = 24'h000000;
assign target_only_stripe[6584] = 24'h000000;
assign target_only_stripe[6585] = 24'h000000;
assign target_only_stripe[6586] = 24'h000000;
assign target_only_stripe[6587] = 24'h000000;
assign target_only_stripe[6588] = 24'h000000;
assign target_only_stripe[6589] = 24'h000000;
assign target_only_stripe[6590] = 24'h000000;
assign target_only_stripe[6591] = 24'h000000;
assign target_only_stripe[6592] = 24'h000000;
assign target_only_stripe[6593] = 24'h000000;
assign target_only_stripe[6594] = 24'h000000;
assign target_only_stripe[6595] = 24'h000000;
assign target_only_stripe[6596] = 24'h000000;
assign target_only_stripe[6597] = 24'h000000;
assign target_only_stripe[6598] = 24'h000000;
assign target_only_stripe[6599] = 24'h000000;
assign target_only_stripe[6600] = 24'h000000;
assign target_only_stripe[6601] = 24'h000000;
assign target_only_stripe[6602] = 24'h000000;
assign target_only_stripe[6603] = 24'h000000;
assign target_only_stripe[6604] = 24'h000000;
assign target_only_stripe[6605] = 24'h000000;
assign target_only_stripe[6606] = 24'h000000;
assign target_only_stripe[6607] = 24'h000000;
assign target_only_stripe[6608] = 24'h000000;
assign target_only_stripe[6609] = 24'h000000;
assign target_only_stripe[6610] = 24'h000000;
assign target_only_stripe[6611] = 24'h000000;
assign target_only_stripe[6612] = 24'hbababa;
assign target_only_stripe[6613] = 24'hffffff;
assign target_only_stripe[6614] = 24'hffffff;
assign target_only_stripe[6615] = 24'hffffff;
assign target_only_stripe[6616] = 24'hffffff;
assign target_only_stripe[6617] = 24'hffffff;
assign target_only_stripe[6618] = 24'hffffff;
assign target_only_stripe[6619] = 24'hffffff;
assign target_only_stripe[6620] = 24'hffffff;
assign target_only_stripe[6621] = 24'hffffff;
assign target_only_stripe[6622] = 24'hffffff;
assign target_only_stripe[6623] = 24'hffffff;
assign target_only_stripe[6624] = 24'hffffff;
assign target_only_stripe[6625] = 24'hffffff;
assign target_only_stripe[6626] = 24'hffffff;
assign target_only_stripe[6627] = 24'hffffff;
assign target_only_stripe[6628] = 24'hffffff;
assign target_only_stripe[6629] = 24'hffffff;
assign target_only_stripe[6630] = 24'hffffff;
assign target_only_stripe[6631] = 24'hffffff;
assign target_only_stripe[6632] = 24'hffffff;
assign target_only_stripe[6633] = 24'hffffff;
assign target_only_stripe[6634] = 24'hffffff;
assign target_only_stripe[6635] = 24'hffffff;
assign target_only_stripe[6636] = 24'hffffff;
assign target_only_stripe[6637] = 24'hffffff;
assign target_only_stripe[6638] = 24'hffffff;
assign target_only_stripe[6639] = 24'hffffff;
assign target_only_stripe[6640] = 24'hffffff;
assign target_only_stripe[6641] = 24'hffffff;
assign target_only_stripe[6642] = 24'hffffff;
assign target_only_stripe[6643] = 24'hffffff;
assign target_only_stripe[6644] = 24'hffffff;
assign target_only_stripe[6645] = 24'he9e9e9;
assign target_only_stripe[6646] = 24'h242424;
assign target_only_stripe[6647] = 24'h000000;
assign target_only_stripe[6648] = 24'h000000;
assign target_only_stripe[6649] = 24'h000000;
assign target_only_stripe[6650] = 24'h000000;
assign target_only_stripe[6651] = 24'h000000;
assign target_only_stripe[6652] = 24'h000000;
assign target_only_stripe[6653] = 24'h000000;
assign target_only_stripe[6654] = 24'h000000;
assign target_only_stripe[6655] = 24'h000000;
assign target_only_stripe[6656] = 24'h000000;
assign target_only_stripe[6657] = 24'h000000;
assign target_only_stripe[6658] = 24'h000000;
assign target_only_stripe[6659] = 24'h000000;
assign target_only_stripe[6660] = 24'h000000;
assign target_only_stripe[6661] = 24'h000000;
assign target_only_stripe[6662] = 24'h000000;
assign target_only_stripe[6663] = 24'h000000;
assign target_only_stripe[6664] = 24'h000000;
assign target_only_stripe[6665] = 24'h000000;
assign target_only_stripe[6666] = 24'h000000;
assign target_only_stripe[6667] = 24'h000000;
assign target_only_stripe[6668] = 24'h000000;
assign target_only_stripe[6669] = 24'h000000;
assign target_only_stripe[6670] = 24'h000000;
assign target_only_stripe[6671] = 24'h000000;
assign target_only_stripe[6672] = 24'h000000;
assign target_only_stripe[6673] = 24'h000000;
assign target_only_stripe[6674] = 24'h000000;
assign target_only_stripe[6675] = 24'h000000;
assign target_only_stripe[6676] = 24'h000000;
assign target_only_stripe[6677] = 24'h000000;
assign target_only_stripe[6678] = 24'h202020;
assign target_only_stripe[6679] = 24'hffffff;
assign target_only_stripe[6680] = 24'hffffff;
assign target_only_stripe[6681] = 24'hffffff;
assign target_only_stripe[6682] = 24'hffffff;
assign target_only_stripe[6683] = 24'hffffff;
assign target_only_stripe[6684] = 24'hffffff;
assign target_only_stripe[6685] = 24'hffffff;
assign target_only_stripe[6686] = 24'hffffff;
assign target_only_stripe[6687] = 24'hffffff;
assign target_only_stripe[6688] = 24'hffffff;
assign target_only_stripe[6689] = 24'hffffff;
assign target_only_stripe[6690] = 24'hffffff;
assign target_only_stripe[6691] = 24'hffffff;
assign target_only_stripe[6692] = 24'hffffff;
assign target_only_stripe[6693] = 24'hffffff;
assign target_only_stripe[6694] = 24'hffffff;
assign target_only_stripe[6695] = 24'hffffff;
assign target_only_stripe[6696] = 24'hffffff;
assign target_only_stripe[6697] = 24'hffffff;
assign target_only_stripe[6698] = 24'hffffff;
assign target_only_stripe[6699] = 24'hffffff;
assign target_only_stripe[6700] = 24'hffffff;
assign target_only_stripe[6701] = 24'hffffff;
assign target_only_stripe[6702] = 24'hffffff;
assign target_only_stripe[6703] = 24'hffffff;
assign target_only_stripe[6704] = 24'hffffff;
assign target_only_stripe[6705] = 24'hffffff;
assign target_only_stripe[6706] = 24'hffffff;
assign target_only_stripe[6707] = 24'hffffff;
assign target_only_stripe[6708] = 24'hffffff;
assign target_only_stripe[6709] = 24'hffffff;
assign target_only_stripe[6710] = 24'hffffff;
assign target_only_stripe[6711] = 24'hffffff;
assign target_only_stripe[6712] = 24'hffffff;
assign target_only_stripe[6713] = 24'h939393;
assign target_only_stripe[6714] = 24'h000000;
assign target_only_stripe[6715] = 24'h000000;
assign target_only_stripe[6716] = 24'h000000;
assign target_only_stripe[6717] = 24'h000000;
assign target_only_stripe[6718] = 24'h000000;
assign target_only_stripe[6719] = 24'h000000;
assign target_only_stripe[6720] = 24'h000000;
assign target_only_stripe[6721] = 24'h000000;
assign target_only_stripe[6722] = 24'h000000;
assign target_only_stripe[6723] = 24'h000000;
assign target_only_stripe[6724] = 24'h000000;
assign target_only_stripe[6725] = 24'h000000;
assign target_only_stripe[6726] = 24'h000000;
assign target_only_stripe[6727] = 24'h000000;
assign target_only_stripe[6728] = 24'h000000;
assign target_only_stripe[6729] = 24'h000000;
assign target_only_stripe[6730] = 24'h000000;
assign target_only_stripe[6731] = 24'h000000;
assign target_only_stripe[6732] = 24'h000000;
assign target_only_stripe[6733] = 24'h000000;
assign target_only_stripe[6734] = 24'h000000;
assign target_only_stripe[6735] = 24'h000000;
assign target_only_stripe[6736] = 24'h000000;
assign target_only_stripe[6737] = 24'h000000;
assign target_only_stripe[6738] = 24'h000000;
assign target_only_stripe[6739] = 24'h000000;
assign target_only_stripe[6740] = 24'h000000;
assign target_only_stripe[6741] = 24'h000000;
assign target_only_stripe[6742] = 24'h000000;
assign target_only_stripe[6743] = 24'h000000;
assign target_only_stripe[6744] = 24'h000000;
assign target_only_stripe[6745] = 24'h000000;
assign target_only_stripe[6746] = 24'h000000;
assign target_only_stripe[6747] = 24'h000000;
assign target_only_stripe[6748] = 24'h000000;
assign target_only_stripe[6749] = 24'h000000;
assign target_only_stripe[6750] = 24'h000000;
assign target_only_stripe[6751] = 24'h000000;
assign target_only_stripe[6752] = 24'h000000;
assign target_only_stripe[6753] = 24'h000000;
assign target_only_stripe[6754] = 24'h000000;
assign target_only_stripe[6755] = 24'h000000;
assign target_only_stripe[6756] = 24'h000000;
assign target_only_stripe[6757] = 24'h000000;
assign target_only_stripe[6758] = 24'h000000;
assign target_only_stripe[6759] = 24'h000000;
assign target_only_stripe[6760] = 24'h000000;
assign target_only_stripe[6761] = 24'h000000;
assign target_only_stripe[6762] = 24'h000000;
assign target_only_stripe[6763] = 24'h000000;
assign target_only_stripe[6764] = 24'h000000;
assign target_only_stripe[6765] = 24'h000000;
assign target_only_stripe[6766] = 24'h000000;
assign target_only_stripe[6767] = 24'h000000;
assign target_only_stripe[6768] = 24'h000000;
assign target_only_stripe[6769] = 24'h000000;
assign target_only_stripe[6770] = 24'h000000;
assign target_only_stripe[6771] = 24'h000000;
assign target_only_stripe[6772] = 24'h000000;
assign target_only_stripe[6773] = 24'h000000;
assign target_only_stripe[6774] = 24'h000000;
assign target_only_stripe[6775] = 24'h8b8b8b;
assign target_only_stripe[6776] = 24'hffffff;
assign target_only_stripe[6777] = 24'hffffff;
assign target_only_stripe[6778] = 24'hffffff;
assign target_only_stripe[6779] = 24'hffffff;
assign target_only_stripe[6780] = 24'hffffff;
assign target_only_stripe[6781] = 24'hffffff;
assign target_only_stripe[6782] = 24'hffffff;
assign target_only_stripe[6783] = 24'hffffff;
assign target_only_stripe[6784] = 24'hffffff;
assign target_only_stripe[6785] = 24'hffffff;
assign target_only_stripe[6786] = 24'hffffff;
assign target_only_stripe[6787] = 24'hffffff;
assign target_only_stripe[6788] = 24'hffffff;
assign target_only_stripe[6789] = 24'hffffff;
assign target_only_stripe[6790] = 24'hffffff;
assign target_only_stripe[6791] = 24'hffffff;
assign target_only_stripe[6792] = 24'hffffff;
assign target_only_stripe[6793] = 24'hffffff;
assign target_only_stripe[6794] = 24'hffffff;
assign target_only_stripe[6795] = 24'hffffff;
assign target_only_stripe[6796] = 24'hffffff;
assign target_only_stripe[6797] = 24'hffffff;
assign target_only_stripe[6798] = 24'hffffff;
assign target_only_stripe[6799] = 24'hffffff;
assign target_only_stripe[6800] = 24'hffffff;
assign target_only_stripe[6801] = 24'hffffff;
assign target_only_stripe[6802] = 24'hffffff;
assign target_only_stripe[6803] = 24'hffffff;
assign target_only_stripe[6804] = 24'hffffff;
assign target_only_stripe[6805] = 24'hffffff;
assign target_only_stripe[6806] = 24'hffffff;
assign target_only_stripe[6807] = 24'hffffff;
assign target_only_stripe[6808] = 24'hffffff;
assign target_only_stripe[6809] = 24'hffffff;
assign target_only_stripe[6810] = 24'h262626;
assign target_only_stripe[6811] = 24'h000000;
assign target_only_stripe[6812] = 24'h000000;
assign target_only_stripe[6813] = 24'h000000;
assign target_only_stripe[6814] = 24'h000000;
assign target_only_stripe[6815] = 24'h000000;
assign target_only_stripe[6816] = 24'h000000;
assign target_only_stripe[6817] = 24'h000000;
assign target_only_stripe[6818] = 24'h000000;
assign target_only_stripe[6819] = 24'h000000;
assign target_only_stripe[6820] = 24'h000000;
assign target_only_stripe[6821] = 24'h000000;
assign target_only_stripe[6822] = 24'h000000;
assign target_only_stripe[6823] = 24'h000000;
assign target_only_stripe[6824] = 24'h000000;
assign target_only_stripe[6825] = 24'h000000;
assign target_only_stripe[6826] = 24'h000000;
assign target_only_stripe[6827] = 24'h000000;
assign target_only_stripe[6828] = 24'h000000;
assign target_only_stripe[6829] = 24'h000000;
assign target_only_stripe[6830] = 24'h000000;
assign target_only_stripe[6831] = 24'h000000;
assign target_only_stripe[6832] = 24'h000000;
assign target_only_stripe[6833] = 24'h000000;
assign target_only_stripe[6834] = 24'h000000;
assign target_only_stripe[6835] = 24'h000000;
assign target_only_stripe[6836] = 24'h000000;
assign target_only_stripe[6837] = 24'h000000;
assign target_only_stripe[6838] = 24'h000000;
assign target_only_stripe[6839] = 24'h000000;
assign target_only_stripe[6840] = 24'h000000;
assign target_only_stripe[6841] = 24'h000000;
assign target_only_stripe[6842] = 24'h1b1b1b;
assign target_only_stripe[6843] = 24'he5e5e5;
assign target_only_stripe[6844] = 24'hffffff;
assign target_only_stripe[6845] = 24'hffffff;
assign target_only_stripe[6846] = 24'hffffff;
assign target_only_stripe[6847] = 24'hffffff;
assign target_only_stripe[6848] = 24'hffffff;
assign target_only_stripe[6849] = 24'hffffff;
assign target_only_stripe[6850] = 24'hffffff;
assign target_only_stripe[6851] = 24'hffffff;
assign target_only_stripe[6852] = 24'hffffff;
assign target_only_stripe[6853] = 24'hffffff;
assign target_only_stripe[6854] = 24'hffffff;
assign target_only_stripe[6855] = 24'hffffff;
assign target_only_stripe[6856] = 24'hffffff;
assign target_only_stripe[6857] = 24'hffffff;
assign target_only_stripe[6858] = 24'hffffff;
assign target_only_stripe[6859] = 24'hffffff;
assign target_only_stripe[6860] = 24'hffffff;
assign target_only_stripe[6861] = 24'hffffff;
assign target_only_stripe[6862] = 24'hffffff;
assign target_only_stripe[6863] = 24'hffffff;
assign target_only_stripe[6864] = 24'hffffff;
assign target_only_stripe[6865] = 24'hffffff;
assign target_only_stripe[6866] = 24'hffffff;
assign target_only_stripe[6867] = 24'hffffff;
assign target_only_stripe[6868] = 24'hffffff;
assign target_only_stripe[6869] = 24'hffffff;
assign target_only_stripe[6870] = 24'hfaf7f5;
assign target_only_stripe[6871] = 24'hffffff;
assign target_only_stripe[6872] = 24'hffffff;
assign target_only_stripe[6873] = 24'hffffff;
assign target_only_stripe[6874] = 24'hffffff;
assign target_only_stripe[6875] = 24'hffffff;
assign target_only_stripe[6876] = 24'hc0c0c0;
assign target_only_stripe[6877] = 24'h000000;
assign target_only_stripe[6878] = 24'h000000;
assign target_only_stripe[6879] = 24'h000000;
assign target_only_stripe[6880] = 24'h000000;
assign target_only_stripe[6881] = 24'h000000;
assign target_only_stripe[6882] = 24'h000000;
assign target_only_stripe[6883] = 24'h000000;
assign target_only_stripe[6884] = 24'h000000;
assign target_only_stripe[6885] = 24'h000000;
assign target_only_stripe[6886] = 24'h000000;
assign target_only_stripe[6887] = 24'h000000;
assign target_only_stripe[6888] = 24'h000000;
assign target_only_stripe[6889] = 24'h000000;
assign target_only_stripe[6890] = 24'h000000;
assign target_only_stripe[6891] = 24'h000000;
assign target_only_stripe[6892] = 24'h000000;
assign target_only_stripe[6893] = 24'h000000;
assign target_only_stripe[6894] = 24'h000000;
assign target_only_stripe[6895] = 24'h000000;
assign target_only_stripe[6896] = 24'h000000;
assign target_only_stripe[6897] = 24'h000000;
assign target_only_stripe[6898] = 24'h000000;
assign target_only_stripe[6899] = 24'h000000;
assign target_only_stripe[6900] = 24'h000000;
assign target_only_stripe[6901] = 24'h000000;
assign target_only_stripe[6902] = 24'h000000;
assign target_only_stripe[6903] = 24'h000000;
assign target_only_stripe[6904] = 24'h000000;
assign target_only_stripe[6905] = 24'h000000;
assign target_only_stripe[6906] = 24'h000000;
assign target_only_stripe[6907] = 24'h000000;
assign target_only_stripe[6908] = 24'h000000;
assign target_only_stripe[6909] = 24'h000000;
assign target_only_stripe[6910] = 24'h000000;
assign target_only_stripe[6911] = 24'h000000;
assign target_only_stripe[6912] = 24'h000000;
assign target_only_stripe[6913] = 24'h000000;
assign target_only_stripe[6914] = 24'h000000;
assign target_only_stripe[6915] = 24'h000000;
assign target_only_stripe[6916] = 24'h000000;
assign target_only_stripe[6917] = 24'h000000;
assign target_only_stripe[6918] = 24'h000000;
assign target_only_stripe[6919] = 24'h000000;
assign target_only_stripe[6920] = 24'h000000;
assign target_only_stripe[6921] = 24'h000000;
assign target_only_stripe[6922] = 24'h000000;
assign target_only_stripe[6923] = 24'h000000;
assign target_only_stripe[6924] = 24'h000000;
assign target_only_stripe[6925] = 24'h000000;
assign target_only_stripe[6926] = 24'h000000;
assign target_only_stripe[6927] = 24'h000000;
assign target_only_stripe[6928] = 24'h000000;
assign target_only_stripe[6929] = 24'h000000;
assign target_only_stripe[6930] = 24'h000000;
assign target_only_stripe[6931] = 24'h000000;
assign target_only_stripe[6932] = 24'h000000;
assign target_only_stripe[6933] = 24'h000000;
assign target_only_stripe[6934] = 24'h000000;
assign target_only_stripe[6935] = 24'h000000;
assign target_only_stripe[6936] = 24'h000000;
assign target_only_stripe[6937] = 24'h000000;
assign target_only_stripe[6938] = 24'h000000;
assign target_only_stripe[6939] = 24'h000000;
assign target_only_stripe[6940] = 24'h000000;
assign target_only_stripe[6941] = 24'hb4b4b4;
assign target_only_stripe[6942] = 24'hffffff;
assign target_only_stripe[6943] = 24'hffffff;
assign target_only_stripe[6944] = 24'hffffff;
assign target_only_stripe[6945] = 24'hffffff;
assign target_only_stripe[6946] = 24'hffffff;
assign target_only_stripe[6947] = 24'hffffff;
assign target_only_stripe[6948] = 24'hffffff;
assign target_only_stripe[6949] = 24'hffffff;
assign target_only_stripe[6950] = 24'hffffff;
assign target_only_stripe[6951] = 24'hffffff;
assign target_only_stripe[6952] = 24'hffffff;
assign target_only_stripe[6953] = 24'hffffff;
assign target_only_stripe[6954] = 24'hffffff;
assign target_only_stripe[6955] = 24'hffffff;
assign target_only_stripe[6956] = 24'hffffff;
assign target_only_stripe[6957] = 24'hffffff;
assign target_only_stripe[6958] = 24'hffffff;
assign target_only_stripe[6959] = 24'hffffff;
assign target_only_stripe[6960] = 24'hffffff;
assign target_only_stripe[6961] = 24'hffffff;
assign target_only_stripe[6962] = 24'hffffff;
assign target_only_stripe[6963] = 24'hffffff;
assign target_only_stripe[6964] = 24'hffffff;
assign target_only_stripe[6965] = 24'hffffff;
assign target_only_stripe[6966] = 24'hffffff;
assign target_only_stripe[6967] = 24'hffffff;
assign target_only_stripe[6968] = 24'hffffff;
assign target_only_stripe[6969] = 24'hffffff;
assign target_only_stripe[6970] = 24'hffffff;
assign target_only_stripe[6971] = 24'hffffff;
assign target_only_stripe[6972] = 24'hffffff;
assign target_only_stripe[6973] = 24'hffffff;
assign target_only_stripe[6974] = 24'hffffff;
assign target_only_stripe[6975] = 24'hd6d6d6;
assign target_only_stripe[6976] = 24'h000000;
assign target_only_stripe[6977] = 24'h000000;
assign target_only_stripe[6978] = 24'h000000;
assign target_only_stripe[6979] = 24'h000000;
assign target_only_stripe[6980] = 24'h000000;
assign target_only_stripe[6981] = 24'h000000;
assign target_only_stripe[6982] = 24'h000000;
assign target_only_stripe[6983] = 24'h000000;
assign target_only_stripe[6984] = 24'h000000;
assign target_only_stripe[6985] = 24'h000000;
assign target_only_stripe[6986] = 24'h000000;
assign target_only_stripe[6987] = 24'h000000;
assign target_only_stripe[6988] = 24'h000000;
assign target_only_stripe[6989] = 24'h000000;
assign target_only_stripe[6990] = 24'h000000;
assign target_only_stripe[6991] = 24'h000000;
assign target_only_stripe[6992] = 24'h000000;
assign target_only_stripe[6993] = 24'h000000;
assign target_only_stripe[6994] = 24'h000000;
assign target_only_stripe[6995] = 24'h000000;
assign target_only_stripe[6996] = 24'h000000;
assign target_only_stripe[6997] = 24'h000000;
assign target_only_stripe[6998] = 24'h000000;
assign target_only_stripe[6999] = 24'h000000;
assign target_only_stripe[7000] = 24'h000000;
assign target_only_stripe[7001] = 24'h000000;
assign target_only_stripe[7002] = 24'h000000;
assign target_only_stripe[7003] = 24'h000000;
assign target_only_stripe[7004] = 24'h000000;
assign target_only_stripe[7005] = 24'h000000;
assign target_only_stripe[7006] = 24'h000000;
assign target_only_stripe[7007] = 24'h030303;
assign target_only_stripe[7008] = 24'hffffff;
assign target_only_stripe[7009] = 24'hffffff;
assign target_only_stripe[7010] = 24'hffffff;
assign target_only_stripe[7011] = 24'hffffff;
assign target_only_stripe[7012] = 24'hffffff;
assign target_only_stripe[7013] = 24'hffffff;
assign target_only_stripe[7014] = 24'hffffff;
assign target_only_stripe[7015] = 24'hffffff;
assign target_only_stripe[7016] = 24'hffffff;
assign target_only_stripe[7017] = 24'hffffff;
assign target_only_stripe[7018] = 24'hffffff;
assign target_only_stripe[7019] = 24'hffffff;
assign target_only_stripe[7020] = 24'hffffff;
assign target_only_stripe[7021] = 24'hffffff;
assign target_only_stripe[7022] = 24'hffffff;
assign target_only_stripe[7023] = 24'hffffff;
assign target_only_stripe[7024] = 24'hffffff;
assign target_only_stripe[7025] = 24'hffffff;
assign target_only_stripe[7026] = 24'hffffff;
assign target_only_stripe[7027] = 24'hffffff;
assign target_only_stripe[7028] = 24'hffffff;
assign target_only_stripe[7029] = 24'hffffff;
assign target_only_stripe[7030] = 24'hffffff;
assign target_only_stripe[7031] = 24'hffffff;
assign target_only_stripe[7032] = 24'hffffff;
assign target_only_stripe[7033] = 24'hffffff;
assign target_only_stripe[7034] = 24'hffffff;
assign target_only_stripe[7035] = 24'hffffff;
assign target_only_stripe[7036] = 24'hffffff;
assign target_only_stripe[7037] = 24'hffffff;
assign target_only_stripe[7038] = 24'hffffff;
assign target_only_stripe[7039] = 24'hffffff;
assign target_only_stripe[7040] = 24'hffffff;
assign target_only_stripe[7041] = 24'hffffff;
assign target_only_stripe[7042] = 24'hffffff;
assign target_only_stripe[7043] = 24'h090909;
assign target_only_stripe[7044] = 24'h000000;
assign target_only_stripe[7045] = 24'h000000;
assign target_only_stripe[7046] = 24'h000000;
assign target_only_stripe[7047] = 24'h000000;
assign target_only_stripe[7048] = 24'h000000;
assign target_only_stripe[7049] = 24'h000000;
assign target_only_stripe[7050] = 24'h000000;
assign target_only_stripe[7051] = 24'h000000;
assign target_only_stripe[7052] = 24'h000000;
assign target_only_stripe[7053] = 24'h000000;
assign target_only_stripe[7054] = 24'h000000;
assign target_only_stripe[7055] = 24'h000000;
assign target_only_stripe[7056] = 24'h000000;
assign target_only_stripe[7057] = 24'h000000;
assign target_only_stripe[7058] = 24'h000000;
assign target_only_stripe[7059] = 24'h000000;
assign target_only_stripe[7060] = 24'h000000;
assign target_only_stripe[7061] = 24'h000000;
assign target_only_stripe[7062] = 24'h000000;
assign target_only_stripe[7063] = 24'h000000;
assign target_only_stripe[7064] = 24'h000000;
assign target_only_stripe[7065] = 24'h000000;
assign target_only_stripe[7066] = 24'h000000;
assign target_only_stripe[7067] = 24'h000000;
assign target_only_stripe[7068] = 24'h000000;
assign target_only_stripe[7069] = 24'h000000;
assign target_only_stripe[7070] = 24'h000000;
assign target_only_stripe[7071] = 24'h000000;
assign target_only_stripe[7072] = 24'h000000;
assign target_only_stripe[7073] = 24'h000000;
assign target_only_stripe[7074] = 24'h000000;
assign target_only_stripe[7075] = 24'h000000;
assign target_only_stripe[7076] = 24'h000000;
assign target_only_stripe[7077] = 24'h000000;
assign target_only_stripe[7078] = 24'h000000;
assign target_only_stripe[7079] = 24'h000000;
assign target_only_stripe[7080] = 24'h000000;
assign target_only_stripe[7081] = 24'h000000;
assign target_only_stripe[7082] = 24'h000000;
assign target_only_stripe[7083] = 24'h000000;
assign target_only_stripe[7084] = 24'h000000;
assign target_only_stripe[7085] = 24'h000000;
assign target_only_stripe[7086] = 24'h000000;
assign target_only_stripe[7087] = 24'h000000;
assign target_only_stripe[7088] = 24'h000000;
assign target_only_stripe[7089] = 24'h000000;
assign target_only_stripe[7090] = 24'h000000;
assign target_only_stripe[7091] = 24'h000000;
assign target_only_stripe[7092] = 24'h000000;
assign target_only_stripe[7093] = 24'h000000;
assign target_only_stripe[7094] = 24'h000000;
assign target_only_stripe[7095] = 24'h000000;
assign target_only_stripe[7096] = 24'h000000;
assign target_only_stripe[7097] = 24'h000000;
assign target_only_stripe[7098] = 24'h000000;
assign target_only_stripe[7099] = 24'h000000;
assign target_only_stripe[7100] = 24'h000000;
assign target_only_stripe[7101] = 24'h000000;
assign target_only_stripe[7102] = 24'h000000;
assign target_only_stripe[7103] = 24'h060606;
assign target_only_stripe[7104] = 24'hf7f7f7;
assign target_only_stripe[7105] = 24'hffffff;
assign target_only_stripe[7106] = 24'hffffff;
assign target_only_stripe[7107] = 24'hffffff;
assign target_only_stripe[7108] = 24'hffffff;
assign target_only_stripe[7109] = 24'hffffff;
assign target_only_stripe[7110] = 24'hffffff;
assign target_only_stripe[7111] = 24'hffffff;
assign target_only_stripe[7112] = 24'hffffff;
assign target_only_stripe[7113] = 24'hffffff;
assign target_only_stripe[7114] = 24'hffffff;
assign target_only_stripe[7115] = 24'hffffff;
assign target_only_stripe[7116] = 24'hffffff;
assign target_only_stripe[7117] = 24'hffffff;
assign target_only_stripe[7118] = 24'hffffff;
assign target_only_stripe[7119] = 24'hffffff;
assign target_only_stripe[7120] = 24'hffffff;
assign target_only_stripe[7121] = 24'hffffff;
assign target_only_stripe[7122] = 24'hffffff;
assign target_only_stripe[7123] = 24'hffffff;
assign target_only_stripe[7124] = 24'hffffff;
assign target_only_stripe[7125] = 24'hffffff;
assign target_only_stripe[7126] = 24'hffffff;
assign target_only_stripe[7127] = 24'hffffff;
assign target_only_stripe[7128] = 24'hffffff;
assign target_only_stripe[7129] = 24'hffffff;
assign target_only_stripe[7130] = 24'hffffff;
assign target_only_stripe[7131] = 24'hffffff;
assign target_only_stripe[7132] = 24'hffffff;
assign target_only_stripe[7133] = 24'hffffff;
assign target_only_stripe[7134] = 24'hffffff;
assign target_only_stripe[7135] = 24'hffffff;
assign target_only_stripe[7136] = 24'hffffff;
assign target_only_stripe[7137] = 24'hffffff;
assign target_only_stripe[7138] = 24'hffffff;
assign target_only_stripe[7139] = 24'h040404;
assign target_only_stripe[7140] = 24'h000000;
assign target_only_stripe[7141] = 24'h000000;
assign target_only_stripe[7142] = 24'h000000;
assign target_only_stripe[7143] = 24'h000000;
assign target_only_stripe[7144] = 24'h000000;
assign target_only_stripe[7145] = 24'h000000;
assign target_only_stripe[7146] = 24'h000000;
assign target_only_stripe[7147] = 24'h000000;
assign target_only_stripe[7148] = 24'h000000;
assign target_only_stripe[7149] = 24'h000000;
assign target_only_stripe[7150] = 24'h000000;
assign target_only_stripe[7151] = 24'h000000;
assign target_only_stripe[7152] = 24'h000000;
assign target_only_stripe[7153] = 24'h000000;
assign target_only_stripe[7154] = 24'h000000;
assign target_only_stripe[7155] = 24'h000000;
assign target_only_stripe[7156] = 24'h000000;
assign target_only_stripe[7157] = 24'h000000;
assign target_only_stripe[7158] = 24'h000000;
assign target_only_stripe[7159] = 24'h000000;
assign target_only_stripe[7160] = 24'h000000;
assign target_only_stripe[7161] = 24'h000000;
assign target_only_stripe[7162] = 24'h000000;
assign target_only_stripe[7163] = 24'h000000;
assign target_only_stripe[7164] = 24'h000000;
assign target_only_stripe[7165] = 24'h000000;
assign target_only_stripe[7166] = 24'h000000;
assign target_only_stripe[7167] = 24'h000000;
assign target_only_stripe[7168] = 24'h000000;
assign target_only_stripe[7169] = 24'h000000;
assign target_only_stripe[7170] = 24'h000000;
assign target_only_stripe[7171] = 24'hb4b4b4;
assign target_only_stripe[7172] = 24'hffffff;
assign target_only_stripe[7173] = 24'hffffff;
assign target_only_stripe[7174] = 24'hffffff;
assign target_only_stripe[7175] = 24'hffffff;
assign target_only_stripe[7176] = 24'hffffff;
assign target_only_stripe[7177] = 24'hffffff;
assign target_only_stripe[7178] = 24'hffffff;
assign target_only_stripe[7179] = 24'hffffff;
assign target_only_stripe[7180] = 24'hffffff;
assign target_only_stripe[7181] = 24'hffffff;
assign target_only_stripe[7182] = 24'hffffff;
assign target_only_stripe[7183] = 24'hffffff;
assign target_only_stripe[7184] = 24'hffffff;
assign target_only_stripe[7185] = 24'hffffff;
assign target_only_stripe[7186] = 24'hffffff;
assign target_only_stripe[7187] = 24'hffffff;
assign target_only_stripe[7188] = 24'hffffff;
assign target_only_stripe[7189] = 24'hffffff;
assign target_only_stripe[7190] = 24'hffffff;
assign target_only_stripe[7191] = 24'hffffff;
assign target_only_stripe[7192] = 24'hffffff;
assign target_only_stripe[7193] = 24'hffffff;
assign target_only_stripe[7194] = 24'hffffff;
assign target_only_stripe[7195] = 24'hffffff;
assign target_only_stripe[7196] = 24'hffffff;
assign target_only_stripe[7197] = 24'hffffff;
assign target_only_stripe[7198] = 24'hffffff;
assign target_only_stripe[7199] = 24'hffffff;
assign target_only_stripe[7200] = 24'hffffff;
assign target_only_stripe[7201] = 24'hffffff;
assign target_only_stripe[7202] = 24'hffffff;
assign target_only_stripe[7203] = 24'hffffff;
assign target_only_stripe[7204] = 24'hffffff;
assign target_only_stripe[7205] = 24'hbababa;
assign target_only_stripe[7206] = 24'h000000;
assign target_only_stripe[7207] = 24'h000000;
assign target_only_stripe[7208] = 24'h000000;
assign target_only_stripe[7209] = 24'h000000;
assign target_only_stripe[7210] = 24'h000000;
assign target_only_stripe[7211] = 24'h000000;
assign target_only_stripe[7212] = 24'h000000;
assign target_only_stripe[7213] = 24'h000000;
assign target_only_stripe[7214] = 24'h000000;
assign target_only_stripe[7215] = 24'h000000;
assign target_only_stripe[7216] = 24'h000000;
assign target_only_stripe[7217] = 24'h000000;
assign target_only_stripe[7218] = 24'h000000;
assign target_only_stripe[7219] = 24'h000000;
assign target_only_stripe[7220] = 24'h000000;
assign target_only_stripe[7221] = 24'h000000;
assign target_only_stripe[7222] = 24'h000000;
assign target_only_stripe[7223] = 24'h000000;
assign target_only_stripe[7224] = 24'h000000;
assign target_only_stripe[7225] = 24'h000000;
assign target_only_stripe[7226] = 24'h000000;
assign target_only_stripe[7227] = 24'h000000;
assign target_only_stripe[7228] = 24'h000000;
assign target_only_stripe[7229] = 24'h000000;
assign target_only_stripe[7230] = 24'h000000;
assign target_only_stripe[7231] = 24'h000000;
assign target_only_stripe[7232] = 24'h000000;
assign target_only_stripe[7233] = 24'h000000;
assign target_only_stripe[7234] = 24'h000000;
assign target_only_stripe[7235] = 24'h000000;
assign target_only_stripe[7236] = 24'h000000;
assign target_only_stripe[7237] = 24'h000000;
assign target_only_stripe[7238] = 24'h000000;
assign target_only_stripe[7239] = 24'h000000;
assign target_only_stripe[7240] = 24'h000000;
assign target_only_stripe[7241] = 24'h000000;
assign target_only_stripe[7242] = 24'h000000;
assign target_only_stripe[7243] = 24'h000000;
assign target_only_stripe[7244] = 24'h000000;
assign target_only_stripe[7245] = 24'h000000;
assign target_only_stripe[7246] = 24'h000000;
assign target_only_stripe[7247] = 24'h000000;
assign target_only_stripe[7248] = 24'h000000;
assign target_only_stripe[7249] = 24'h000000;
assign target_only_stripe[7250] = 24'h000000;
assign target_only_stripe[7251] = 24'h000000;
assign target_only_stripe[7252] = 24'h000000;
assign target_only_stripe[7253] = 24'h000000;
assign target_only_stripe[7254] = 24'h000000;
assign target_only_stripe[7255] = 24'h000000;
assign target_only_stripe[7256] = 24'h000000;
assign target_only_stripe[7257] = 24'h000000;
assign target_only_stripe[7258] = 24'h000000;
assign target_only_stripe[7259] = 24'h000000;
assign target_only_stripe[7260] = 24'h000000;
assign target_only_stripe[7261] = 24'h000000;
assign target_only_stripe[7262] = 24'h000000;
assign target_only_stripe[7263] = 24'h000000;
assign target_only_stripe[7264] = 24'h000000;
assign target_only_stripe[7265] = 24'h000000;
assign target_only_stripe[7266] = 24'h000000;
assign target_only_stripe[7267] = 24'h000000;
assign target_only_stripe[7268] = 24'h000000;
assign target_only_stripe[7269] = 24'h000000;
assign target_only_stripe[7270] = 24'ha8a8a8;
assign target_only_stripe[7271] = 24'hffffff;
assign target_only_stripe[7272] = 24'hffffff;
assign target_only_stripe[7273] = 24'hffffff;
assign target_only_stripe[7274] = 24'hffffff;
assign target_only_stripe[7275] = 24'hffffff;
assign target_only_stripe[7276] = 24'hffffff;
assign target_only_stripe[7277] = 24'hffffff;
assign target_only_stripe[7278] = 24'hffffff;
assign target_only_stripe[7279] = 24'hffffff;
assign target_only_stripe[7280] = 24'hffffff;
assign target_only_stripe[7281] = 24'hffffff;
assign target_only_stripe[7282] = 24'hffffff;
assign target_only_stripe[7283] = 24'hffffff;
assign target_only_stripe[7284] = 24'hffffff;
assign target_only_stripe[7285] = 24'hffffff;
assign target_only_stripe[7286] = 24'hffffff;
assign target_only_stripe[7287] = 24'hffffff;
assign target_only_stripe[7288] = 24'hffffff;
assign target_only_stripe[7289] = 24'hffffff;
assign target_only_stripe[7290] = 24'hffffff;
assign target_only_stripe[7291] = 24'hffffff;
assign target_only_stripe[7292] = 24'hffffff;
assign target_only_stripe[7293] = 24'hffffff;
assign target_only_stripe[7294] = 24'hffffff;
assign target_only_stripe[7295] = 24'hffffff;
assign target_only_stripe[7296] = 24'hffffff;
assign target_only_stripe[7297] = 24'hffffff;
assign target_only_stripe[7298] = 24'hffffff;
assign target_only_stripe[7299] = 24'hffffff;
assign target_only_stripe[7300] = 24'hffffff;
assign target_only_stripe[7301] = 24'hffffff;
assign target_only_stripe[7302] = 24'hffffff;
assign target_only_stripe[7303] = 24'hffffff;
assign target_only_stripe[7304] = 24'hffffff;
assign target_only_stripe[7305] = 24'h000000;
assign target_only_stripe[7306] = 24'h000000;
assign target_only_stripe[7307] = 24'h000000;
assign target_only_stripe[7308] = 24'h000000;
assign target_only_stripe[7309] = 24'h000000;
assign target_only_stripe[7310] = 24'h000000;
assign target_only_stripe[7311] = 24'h000000;
assign target_only_stripe[7312] = 24'h000000;
assign target_only_stripe[7313] = 24'h000000;
assign target_only_stripe[7314] = 24'h000000;
assign target_only_stripe[7315] = 24'h000000;
assign target_only_stripe[7316] = 24'h000000;
assign target_only_stripe[7317] = 24'h000000;
assign target_only_stripe[7318] = 24'h000000;
assign target_only_stripe[7319] = 24'h000000;
assign target_only_stripe[7320] = 24'h000000;
assign target_only_stripe[7321] = 24'h000000;
assign target_only_stripe[7322] = 24'h000000;
assign target_only_stripe[7323] = 24'h000000;
assign target_only_stripe[7324] = 24'h000000;
assign target_only_stripe[7325] = 24'h000000;
assign target_only_stripe[7326] = 24'h000000;
assign target_only_stripe[7327] = 24'h000000;
assign target_only_stripe[7328] = 24'h000000;
assign target_only_stripe[7329] = 24'h000000;
assign target_only_stripe[7330] = 24'h000000;
assign target_only_stripe[7331] = 24'h000000;
assign target_only_stripe[7332] = 24'h000000;
assign target_only_stripe[7333] = 24'h000000;
assign target_only_stripe[7334] = 24'h000000;
assign target_only_stripe[7335] = 24'h000000;
assign target_only_stripe[7336] = 24'h000000;
assign target_only_stripe[7337] = 24'hb4b4b4;
assign target_only_stripe[7338] = 24'hffffff;
assign target_only_stripe[7339] = 24'hffffff;
assign target_only_stripe[7340] = 24'hffffff;
assign target_only_stripe[7341] = 24'hffffff;
assign target_only_stripe[7342] = 24'hffffff;
assign target_only_stripe[7343] = 24'hffffff;
assign target_only_stripe[7344] = 24'hffffff;
assign target_only_stripe[7345] = 24'hffffff;
assign target_only_stripe[7346] = 24'hffffff;
assign target_only_stripe[7347] = 24'hffffff;
assign target_only_stripe[7348] = 24'hffffff;
assign target_only_stripe[7349] = 24'hffffff;
assign target_only_stripe[7350] = 24'hffffff;
assign target_only_stripe[7351] = 24'hffffff;
assign target_only_stripe[7352] = 24'hffffff;
assign target_only_stripe[7353] = 24'hffffff;
assign target_only_stripe[7354] = 24'hffffff;
assign target_only_stripe[7355] = 24'hffffff;
assign target_only_stripe[7356] = 24'hffffff;
assign target_only_stripe[7357] = 24'hffffff;
assign target_only_stripe[7358] = 24'hffffff;
assign target_only_stripe[7359] = 24'hffffff;
assign target_only_stripe[7360] = 24'hffffff;
assign target_only_stripe[7361] = 24'hffffff;
assign target_only_stripe[7362] = 24'hffffff;
assign target_only_stripe[7363] = 24'hffffff;
assign target_only_stripe[7364] = 24'hffffff;
assign target_only_stripe[7365] = 24'hffffff;
assign target_only_stripe[7366] = 24'hffffff;
assign target_only_stripe[7367] = 24'hffffff;
assign target_only_stripe[7368] = 24'hffffff;
assign target_only_stripe[7369] = 24'hffffff;
assign target_only_stripe[7370] = 24'hffffff;
assign target_only_stripe[7371] = 24'hffffff;
assign target_only_stripe[7372] = 24'h494949;
assign target_only_stripe[7373] = 24'h000000;
assign target_only_stripe[7374] = 24'h000000;
assign target_only_stripe[7375] = 24'h000000;
assign target_only_stripe[7376] = 24'h000000;
assign target_only_stripe[7377] = 24'h000000;
assign target_only_stripe[7378] = 24'h000000;
assign target_only_stripe[7379] = 24'h000000;
assign target_only_stripe[7380] = 24'h000000;
assign target_only_stripe[7381] = 24'h000000;
assign target_only_stripe[7382] = 24'h000000;
assign target_only_stripe[7383] = 24'h000000;
assign target_only_stripe[7384] = 24'h000000;
assign target_only_stripe[7385] = 24'h000000;
assign target_only_stripe[7386] = 24'h000000;
assign target_only_stripe[7387] = 24'h000000;
assign target_only_stripe[7388] = 24'h000000;
assign target_only_stripe[7389] = 24'h000000;
assign target_only_stripe[7390] = 24'h000000;
assign target_only_stripe[7391] = 24'h000000;
assign target_only_stripe[7392] = 24'h000000;
assign target_only_stripe[7393] = 24'h000000;
assign target_only_stripe[7394] = 24'h000000;
assign target_only_stripe[7395] = 24'h000000;
assign target_only_stripe[7396] = 24'h000000;
assign target_only_stripe[7397] = 24'h000000;
assign target_only_stripe[7398] = 24'h000000;
assign target_only_stripe[7399] = 24'h000000;
assign target_only_stripe[7400] = 24'h000000;
assign target_only_stripe[7401] = 24'h000000;
assign target_only_stripe[7402] = 24'h000000;
assign target_only_stripe[7403] = 24'h000000;
assign target_only_stripe[7404] = 24'h000000;
assign target_only_stripe[7405] = 24'h000000;
assign target_only_stripe[7406] = 24'h000000;
assign target_only_stripe[7407] = 24'h000000;
assign target_only_stripe[7408] = 24'h000000;
assign target_only_stripe[7409] = 24'h000000;
assign target_only_stripe[7410] = 24'h000000;
assign target_only_stripe[7411] = 24'h000000;
assign target_only_stripe[7412] = 24'h000000;
assign target_only_stripe[7413] = 24'h000000;
assign target_only_stripe[7414] = 24'h000000;
assign target_only_stripe[7415] = 24'h000000;
assign target_only_stripe[7416] = 24'h000000;
assign target_only_stripe[7417] = 24'h000000;
assign target_only_stripe[7418] = 24'h000000;
assign target_only_stripe[7419] = 24'h000000;
assign target_only_stripe[7420] = 24'h000000;
assign target_only_stripe[7421] = 24'h000000;
assign target_only_stripe[7422] = 24'h000000;
assign target_only_stripe[7423] = 24'h000000;
assign target_only_stripe[7424] = 24'h000000;
assign target_only_stripe[7425] = 24'h000000;
assign target_only_stripe[7426] = 24'h000000;
assign target_only_stripe[7427] = 24'h000000;
assign target_only_stripe[7428] = 24'h000000;
assign target_only_stripe[7429] = 24'h000000;
assign target_only_stripe[7430] = 24'h000000;
assign target_only_stripe[7431] = 24'h000000;
assign target_only_stripe[7432] = 24'h414141;
assign target_only_stripe[7433] = 24'hd1b6ac;
assign target_only_stripe[7434] = 24'hffffff;
assign target_only_stripe[7435] = 24'hffffff;
assign target_only_stripe[7436] = 24'hffffff;
assign target_only_stripe[7437] = 24'hffffff;
assign target_only_stripe[7438] = 24'hffffff;
assign target_only_stripe[7439] = 24'hffffff;
assign target_only_stripe[7440] = 24'hffffff;
assign target_only_stripe[7441] = 24'hffffff;
assign target_only_stripe[7442] = 24'hffffff;
assign target_only_stripe[7443] = 24'hffffff;
assign target_only_stripe[7444] = 24'hffffff;
assign target_only_stripe[7445] = 24'hffffff;
assign target_only_stripe[7446] = 24'hffffff;
assign target_only_stripe[7447] = 24'hffffff;
assign target_only_stripe[7448] = 24'hffffff;
assign target_only_stripe[7449] = 24'hffffff;
assign target_only_stripe[7450] = 24'hffffff;
assign target_only_stripe[7451] = 24'hffffff;
assign target_only_stripe[7452] = 24'hffffff;
assign target_only_stripe[7453] = 24'hffffff;
assign target_only_stripe[7454] = 24'hffffff;
assign target_only_stripe[7455] = 24'hffffff;
assign target_only_stripe[7456] = 24'hffffff;
assign target_only_stripe[7457] = 24'hffffff;
assign target_only_stripe[7458] = 24'hffffff;
assign target_only_stripe[7459] = 24'hffffff;
assign target_only_stripe[7460] = 24'hffffff;
assign target_only_stripe[7461] = 24'hffffff;
assign target_only_stripe[7462] = 24'hffffff;
assign target_only_stripe[7463] = 24'hffffff;
assign target_only_stripe[7464] = 24'hffffff;
assign target_only_stripe[7465] = 24'hffffff;
assign target_only_stripe[7466] = 24'hffffff;
assign target_only_stripe[7467] = 24'hcdcdcd;
assign target_only_stripe[7468] = 24'h000000;
assign target_only_stripe[7469] = 24'h000000;
assign target_only_stripe[7470] = 24'h000000;
assign target_only_stripe[7471] = 24'h000000;
assign target_only_stripe[7472] = 24'h000000;
assign target_only_stripe[7473] = 24'h000000;
assign target_only_stripe[7474] = 24'h000000;
assign target_only_stripe[7475] = 24'h000000;
assign target_only_stripe[7476] = 24'h000000;
assign target_only_stripe[7477] = 24'h000000;
assign target_only_stripe[7478] = 24'h000000;
assign target_only_stripe[7479] = 24'h000000;
assign target_only_stripe[7480] = 24'h000000;
assign target_only_stripe[7481] = 24'h000000;
assign target_only_stripe[7482] = 24'h000000;
assign target_only_stripe[7483] = 24'h000000;
assign target_only_stripe[7484] = 24'h000000;
assign target_only_stripe[7485] = 24'h000000;
assign target_only_stripe[7486] = 24'h000000;
assign target_only_stripe[7487] = 24'h000000;
assign target_only_stripe[7488] = 24'h000000;
assign target_only_stripe[7489] = 24'h000000;
assign target_only_stripe[7490] = 24'h000000;
assign target_only_stripe[7491] = 24'h000000;
assign target_only_stripe[7492] = 24'h000000;
assign target_only_stripe[7493] = 24'h000000;
assign target_only_stripe[7494] = 24'h000000;
assign target_only_stripe[7495] = 24'h000000;
assign target_only_stripe[7496] = 24'h000000;
assign target_only_stripe[7497] = 24'h000000;
assign target_only_stripe[7498] = 24'h000000;
assign target_only_stripe[7499] = 24'h000000;
assign target_only_stripe[7500] = 24'hffffff;
assign target_only_stripe[7501] = 24'hffffff;
assign target_only_stripe[7502] = 24'hffffff;
assign target_only_stripe[7503] = 24'hffffff;
assign target_only_stripe[7504] = 24'hffffff;
assign target_only_stripe[7505] = 24'hffffff;
assign target_only_stripe[7506] = 24'hffffff;
assign target_only_stripe[7507] = 24'hffffff;
assign target_only_stripe[7508] = 24'hffffff;
assign target_only_stripe[7509] = 24'hffffff;
assign target_only_stripe[7510] = 24'hffffff;
assign target_only_stripe[7511] = 24'hffffff;
assign target_only_stripe[7512] = 24'hffffff;
assign target_only_stripe[7513] = 24'hffffff;
assign target_only_stripe[7514] = 24'hffffff;
assign target_only_stripe[7515] = 24'hffffff;
assign target_only_stripe[7516] = 24'hffffff;
assign target_only_stripe[7517] = 24'hffffff;
assign target_only_stripe[7518] = 24'hffffff;
assign target_only_stripe[7519] = 24'hffffff;
assign target_only_stripe[7520] = 24'hffffff;
assign target_only_stripe[7521] = 24'hffffff;
assign target_only_stripe[7522] = 24'hffffff;
assign target_only_stripe[7523] = 24'hffffff;
assign target_only_stripe[7524] = 24'hffffff;
assign target_only_stripe[7525] = 24'hffffff;
assign target_only_stripe[7526] = 24'hffffff;
assign target_only_stripe[7527] = 24'hffffff;
assign target_only_stripe[7528] = 24'hffffff;
assign target_only_stripe[7529] = 24'hffffff;
assign target_only_stripe[7530] = 24'hffffff;
assign target_only_stripe[7531] = 24'hffffff;
assign target_only_stripe[7532] = 24'hffffff;
assign target_only_stripe[7533] = 24'hffffff;
assign target_only_stripe[7534] = 24'haeaeae;
assign target_only_stripe[7535] = 24'h000000;
assign target_only_stripe[7536] = 24'h000000;
assign target_only_stripe[7537] = 24'h000000;
assign target_only_stripe[7538] = 24'h000000;
assign target_only_stripe[7539] = 24'h000000;
assign target_only_stripe[7540] = 24'h000000;
assign target_only_stripe[7541] = 24'h000000;
assign target_only_stripe[7542] = 24'h000000;
assign target_only_stripe[7543] = 24'h000000;
assign target_only_stripe[7544] = 24'h000000;
assign target_only_stripe[7545] = 24'h000000;
assign target_only_stripe[7546] = 24'h000000;
assign target_only_stripe[7547] = 24'h000000;
assign target_only_stripe[7548] = 24'h000000;
assign target_only_stripe[7549] = 24'h000000;
assign target_only_stripe[7550] = 24'h000000;
assign target_only_stripe[7551] = 24'h000000;
assign target_only_stripe[7552] = 24'h000000;
assign target_only_stripe[7553] = 24'h000000;
assign target_only_stripe[7554] = 24'h000000;
assign target_only_stripe[7555] = 24'h000000;
assign target_only_stripe[7556] = 24'h000000;
assign target_only_stripe[7557] = 24'h000000;
assign target_only_stripe[7558] = 24'h000000;
assign target_only_stripe[7559] = 24'h000000;
assign target_only_stripe[7560] = 24'h000000;
assign target_only_stripe[7561] = 24'h000000;
assign target_only_stripe[7562] = 24'h000000;
assign target_only_stripe[7563] = 24'h000000;
assign target_only_stripe[7564] = 24'h000000;
assign target_only_stripe[7565] = 24'h000000;
assign target_only_stripe[7566] = 24'h000000;
assign target_only_stripe[7567] = 24'h000000;
assign target_only_stripe[7568] = 24'h000000;
assign target_only_stripe[7569] = 24'h000000;
assign target_only_stripe[7570] = 24'h000000;
assign target_only_stripe[7571] = 24'h000000;
assign target_only_stripe[7572] = 24'h000000;
assign target_only_stripe[7573] = 24'h000000;
assign target_only_stripe[7574] = 24'h000000;
assign target_only_stripe[7575] = 24'h000000;
assign target_only_stripe[7576] = 24'h000000;
assign target_only_stripe[7577] = 24'h000000;
assign target_only_stripe[7578] = 24'h000000;
assign target_only_stripe[7579] = 24'h000000;
assign target_only_stripe[7580] = 24'h000000;
assign target_only_stripe[7581] = 24'h000000;
assign target_only_stripe[7582] = 24'h000000;
assign target_only_stripe[7583] = 24'h000000;
assign target_only_stripe[7584] = 24'h000000;
assign target_only_stripe[7585] = 24'h000000;
assign target_only_stripe[7586] = 24'h000000;
assign target_only_stripe[7587] = 24'h000000;
assign target_only_stripe[7588] = 24'h000000;
assign target_only_stripe[7589] = 24'h000000;
assign target_only_stripe[7590] = 24'h000000;
assign target_only_stripe[7591] = 24'h000000;
assign target_only_stripe[7592] = 24'h000000;
assign target_only_stripe[7593] = 24'h000000;
assign target_only_stripe[7594] = 24'h000000;
assign target_only_stripe[7595] = 24'h000000;
assign target_only_stripe[7596] = 24'h000000;
assign target_only_stripe[7597] = 24'h000000;
assign target_only_stripe[7598] = 24'h000000;
assign target_only_stripe[7599] = 24'hb2b2b2;
assign target_only_stripe[7600] = 24'hffffff;
assign target_only_stripe[7601] = 24'hffffff;
assign target_only_stripe[7602] = 24'hffffff;
assign target_only_stripe[7603] = 24'hffffff;
assign target_only_stripe[7604] = 24'hffffff;
assign target_only_stripe[7605] = 24'hffffff;
assign target_only_stripe[7606] = 24'hffffff;
assign target_only_stripe[7607] = 24'hffffff;
assign target_only_stripe[7608] = 24'hffffff;
assign target_only_stripe[7609] = 24'hffffff;
assign target_only_stripe[7610] = 24'hffffff;
assign target_only_stripe[7611] = 24'hffffff;
assign target_only_stripe[7612] = 24'hffffff;
assign target_only_stripe[7613] = 24'hffffff;
assign target_only_stripe[7614] = 24'hffffff;
assign target_only_stripe[7615] = 24'hffffff;
assign target_only_stripe[7616] = 24'hffffff;
assign target_only_stripe[7617] = 24'hffffff;
assign target_only_stripe[7618] = 24'hffffff;
assign target_only_stripe[7619] = 24'hffffff;
assign target_only_stripe[7620] = 24'hffffff;
assign target_only_stripe[7621] = 24'hffffff;
assign target_only_stripe[7622] = 24'hffffff;
assign target_only_stripe[7623] = 24'hffffff;
assign target_only_stripe[7624] = 24'hffffff;
assign target_only_stripe[7625] = 24'hffffff;
assign target_only_stripe[7626] = 24'hffffff;
assign target_only_stripe[7627] = 24'hffffff;
assign target_only_stripe[7628] = 24'hffffff;
assign target_only_stripe[7629] = 24'hffffff;
assign target_only_stripe[7630] = 24'hffffff;
assign target_only_stripe[7631] = 24'hffffff;
assign target_only_stripe[7632] = 24'hffffff;
assign target_only_stripe[7633] = 24'hffffff;
assign target_only_stripe[7634] = 24'h000000;
assign target_only_stripe[7635] = 24'h000000;
assign target_only_stripe[7636] = 24'h000000;
assign target_only_stripe[7637] = 24'h000000;
assign target_only_stripe[7638] = 24'h000000;
assign target_only_stripe[7639] = 24'h000000;
assign target_only_stripe[7640] = 24'h000000;
assign target_only_stripe[7641] = 24'h000000;
assign target_only_stripe[7642] = 24'h000000;
assign target_only_stripe[7643] = 24'h000000;
assign target_only_stripe[7644] = 24'h000000;
assign target_only_stripe[7645] = 24'h000000;
assign target_only_stripe[7646] = 24'h000000;
assign target_only_stripe[7647] = 24'h000000;
assign target_only_stripe[7648] = 24'h000000;
assign target_only_stripe[7649] = 24'h000000;
assign target_only_stripe[7650] = 24'h000000;
assign target_only_stripe[7651] = 24'h000000;
assign target_only_stripe[7652] = 24'h000000;
assign target_only_stripe[7653] = 24'h000000;
assign target_only_stripe[7654] = 24'h000000;
assign target_only_stripe[7655] = 24'h000000;
assign target_only_stripe[7656] = 24'h000000;
assign target_only_stripe[7657] = 24'h000000;
assign target_only_stripe[7658] = 24'h000000;
assign target_only_stripe[7659] = 24'h000000;
assign target_only_stripe[7660] = 24'h000000;
assign target_only_stripe[7661] = 24'h000000;
assign target_only_stripe[7662] = 24'h000000;
assign target_only_stripe[7663] = 24'h000000;
assign target_only_stripe[7664] = 24'h000000;
assign target_only_stripe[7665] = 24'h000000;
assign target_only_stripe[7666] = 24'h939393;
assign target_only_stripe[7667] = 24'hffffff;
assign target_only_stripe[7668] = 24'hffffff;
assign target_only_stripe[7669] = 24'hffffff;
assign target_only_stripe[7670] = 24'hffffff;
assign target_only_stripe[7671] = 24'hffffff;
assign target_only_stripe[7672] = 24'hffffff;
assign target_only_stripe[7673] = 24'hffffff;
assign target_only_stripe[7674] = 24'hffffff;
assign target_only_stripe[7675] = 24'hffffff;
assign target_only_stripe[7676] = 24'hffffff;
assign target_only_stripe[7677] = 24'hffffff;
assign target_only_stripe[7678] = 24'hffffff;
assign target_only_stripe[7679] = 24'hffffff;
assign target_only_stripe[7680] = 24'hffffff;
assign target_only_stripe[7681] = 24'hffffff;
assign target_only_stripe[7682] = 24'hffffff;
assign target_only_stripe[7683] = 24'hffffff;
assign target_only_stripe[7684] = 24'hffffff;
assign target_only_stripe[7685] = 24'hffffff;
assign target_only_stripe[7686] = 24'hffffff;
assign target_only_stripe[7687] = 24'hffffff;
assign target_only_stripe[7688] = 24'hffffff;
assign target_only_stripe[7689] = 24'hffffff;
assign target_only_stripe[7690] = 24'hffffff;
assign target_only_stripe[7691] = 24'hffffff;
assign target_only_stripe[7692] = 24'hffffff;
assign target_only_stripe[7693] = 24'hffffff;
assign target_only_stripe[7694] = 24'hffffff;
assign target_only_stripe[7695] = 24'hffffff;
assign target_only_stripe[7696] = 24'hffffff;
assign target_only_stripe[7697] = 24'hffffff;
assign target_only_stripe[7698] = 24'hffffff;
assign target_only_stripe[7699] = 24'hffffff;
assign target_only_stripe[7700] = 24'hffffff;
assign target_only_stripe[7701] = 24'h9c9c9c;
assign target_only_stripe[7702] = 24'h000000;
assign target_only_stripe[7703] = 24'h000000;
assign target_only_stripe[7704] = 24'h000000;
assign target_only_stripe[7705] = 24'h000000;
assign target_only_stripe[7706] = 24'h000000;
assign target_only_stripe[7707] = 24'h000000;
assign target_only_stripe[7708] = 24'h000000;
assign target_only_stripe[7709] = 24'h000000;
assign target_only_stripe[7710] = 24'h000000;
assign target_only_stripe[7711] = 24'h000000;
assign target_only_stripe[7712] = 24'h000000;
assign target_only_stripe[7713] = 24'h000000;
assign target_only_stripe[7714] = 24'h000000;
assign target_only_stripe[7715] = 24'h000000;
assign target_only_stripe[7716] = 24'h000000;
assign target_only_stripe[7717] = 24'h000000;
assign target_only_stripe[7718] = 24'h000000;
assign target_only_stripe[7719] = 24'h000000;
assign target_only_stripe[7720] = 24'h000000;
assign target_only_stripe[7721] = 24'h000000;
assign target_only_stripe[7722] = 24'h000000;
assign target_only_stripe[7723] = 24'h000000;
assign target_only_stripe[7724] = 24'h000000;
assign target_only_stripe[7725] = 24'h000000;
assign target_only_stripe[7726] = 24'h000000;
assign target_only_stripe[7727] = 24'h000000;
assign target_only_stripe[7728] = 24'h000000;
assign target_only_stripe[7729] = 24'h000000;
assign target_only_stripe[7730] = 24'h000000;
assign target_only_stripe[7731] = 24'h000000;
assign target_only_stripe[7732] = 24'h000000;
assign target_only_stripe[7733] = 24'h000000;
assign target_only_stripe[7734] = 24'h000000;
assign target_only_stripe[7735] = 24'h000000;
assign target_only_stripe[7736] = 24'h000000;
assign target_only_stripe[7737] = 24'h000000;
assign target_only_stripe[7738] = 24'h000000;
assign target_only_stripe[7739] = 24'h000000;
assign target_only_stripe[7740] = 24'h000000;
assign target_only_stripe[7741] = 24'h000000;
assign target_only_stripe[7742] = 24'h000000;
assign target_only_stripe[7743] = 24'h000000;
assign target_only_stripe[7744] = 24'h000000;
assign target_only_stripe[7745] = 24'h000000;
assign target_only_stripe[7746] = 24'h000000;
assign target_only_stripe[7747] = 24'h000000;
assign target_only_stripe[7748] = 24'h000000;
assign target_only_stripe[7749] = 24'h000000;
assign target_only_stripe[7750] = 24'h000000;
assign target_only_stripe[7751] = 24'h000000;
assign target_only_stripe[7752] = 24'h000000;
assign target_only_stripe[7753] = 24'h000000;
assign target_only_stripe[7754] = 24'h000000;
assign target_only_stripe[7755] = 24'h000000;
assign target_only_stripe[7756] = 24'h000000;
assign target_only_stripe[7757] = 24'h000000;
assign target_only_stripe[7758] = 24'h000000;
assign target_only_stripe[7759] = 24'h000000;
assign target_only_stripe[7760] = 24'h000000;
assign target_only_stripe[7761] = 24'h959595;
assign target_only_stripe[7762] = 24'hffffff;
assign target_only_stripe[7763] = 24'hffffff;
assign target_only_stripe[7764] = 24'hffffff;
assign target_only_stripe[7765] = 24'hffffff;
assign target_only_stripe[7766] = 24'hffffff;
assign target_only_stripe[7767] = 24'hffffff;
assign target_only_stripe[7768] = 24'hffffff;
assign target_only_stripe[7769] = 24'hffffff;
assign target_only_stripe[7770] = 24'hffffff;
assign target_only_stripe[7771] = 24'hffffff;
assign target_only_stripe[7772] = 24'hffffff;
assign target_only_stripe[7773] = 24'hffffff;
assign target_only_stripe[7774] = 24'hffffff;
assign target_only_stripe[7775] = 24'hffffff;
assign target_only_stripe[7776] = 24'hffffff;
assign target_only_stripe[7777] = 24'hffffff;
assign target_only_stripe[7778] = 24'hffffff;
assign target_only_stripe[7779] = 24'hffffff;
assign target_only_stripe[7780] = 24'hffffff;
assign target_only_stripe[7781] = 24'hffffff;
assign target_only_stripe[7782] = 24'hffffff;
assign target_only_stripe[7783] = 24'hffffff;
assign target_only_stripe[7784] = 24'hffffff;
assign target_only_stripe[7785] = 24'hffffff;
assign target_only_stripe[7786] = 24'hffffff;
assign target_only_stripe[7787] = 24'hffffff;
assign target_only_stripe[7788] = 24'hffffff;
assign target_only_stripe[7789] = 24'hffffff;
assign target_only_stripe[7790] = 24'hffffff;
assign target_only_stripe[7791] = 24'hffffff;
assign target_only_stripe[7792] = 24'hffffff;
assign target_only_stripe[7793] = 24'hffffff;
assign target_only_stripe[7794] = 24'hffffff;
assign target_only_stripe[7795] = 24'hffffff;
assign target_only_stripe[7796] = 24'h9b9b9b;
assign target_only_stripe[7797] = 24'h000000;
assign target_only_stripe[7798] = 24'h000000;
assign target_only_stripe[7799] = 24'h000000;
assign target_only_stripe[7800] = 24'h000000;
assign target_only_stripe[7801] = 24'h000000;
assign target_only_stripe[7802] = 24'h000000;
assign target_only_stripe[7803] = 24'h000000;
assign target_only_stripe[7804] = 24'h000000;
assign target_only_stripe[7805] = 24'h000000;
assign target_only_stripe[7806] = 24'h000000;
assign target_only_stripe[7807] = 24'h000000;
assign target_only_stripe[7808] = 24'h000000;
assign target_only_stripe[7809] = 24'h000000;
assign target_only_stripe[7810] = 24'h000000;
assign target_only_stripe[7811] = 24'h000000;
assign target_only_stripe[7812] = 24'h000000;
assign target_only_stripe[7813] = 24'h000000;
assign target_only_stripe[7814] = 24'h000000;
assign target_only_stripe[7815] = 24'h000000;
assign target_only_stripe[7816] = 24'h000000;
assign target_only_stripe[7817] = 24'h000000;
assign target_only_stripe[7818] = 24'h000000;
assign target_only_stripe[7819] = 24'h000000;
assign target_only_stripe[7820] = 24'h000000;
assign target_only_stripe[7821] = 24'h000000;
assign target_only_stripe[7822] = 24'h000000;
assign target_only_stripe[7823] = 24'h000000;
assign target_only_stripe[7824] = 24'h000000;
assign target_only_stripe[7825] = 24'h000000;
assign target_only_stripe[7826] = 24'h000000;
assign target_only_stripe[7827] = 24'h000000;
assign target_only_stripe[7828] = 24'h000000;
assign target_only_stripe[7829] = 24'hffffff;
assign target_only_stripe[7830] = 24'hffffff;
assign target_only_stripe[7831] = 24'hffffff;
assign target_only_stripe[7832] = 24'hffffff;
assign target_only_stripe[7833] = 24'hffffff;
assign target_only_stripe[7834] = 24'hffffff;
assign target_only_stripe[7835] = 24'hffffff;
assign target_only_stripe[7836] = 24'hffffff;
assign target_only_stripe[7837] = 24'hffffff;
assign target_only_stripe[7838] = 24'hffffff;
assign target_only_stripe[7839] = 24'hffffff;
assign target_only_stripe[7840] = 24'hffffff;
assign target_only_stripe[7841] = 24'hffffff;
assign target_only_stripe[7842] = 24'hffffff;
assign target_only_stripe[7843] = 24'hffffff;
assign target_only_stripe[7844] = 24'hffffff;
assign target_only_stripe[7845] = 24'hffffff;
assign target_only_stripe[7846] = 24'hffffff;
assign target_only_stripe[7847] = 24'hffffff;
assign target_only_stripe[7848] = 24'hffffff;
assign target_only_stripe[7849] = 24'hffffff;
assign target_only_stripe[7850] = 24'hffffff;
assign target_only_stripe[7851] = 24'hffffff;
assign target_only_stripe[7852] = 24'hffffff;
assign target_only_stripe[7853] = 24'hffffff;
assign target_only_stripe[7854] = 24'hffffff;
assign target_only_stripe[7855] = 24'hffffff;
assign target_only_stripe[7856] = 24'hffffff;
assign target_only_stripe[7857] = 24'hffffff;
assign target_only_stripe[7858] = 24'hffffff;
assign target_only_stripe[7859] = 24'hffffff;
assign target_only_stripe[7860] = 24'hffffff;
assign target_only_stripe[7861] = 24'hffffff;
assign target_only_stripe[7862] = 24'hffffff;
assign target_only_stripe[7863] = 24'h9c9c9c;
assign target_only_stripe[7864] = 24'h000000;
assign target_only_stripe[7865] = 24'h000000;
assign target_only_stripe[7866] = 24'h000000;
assign target_only_stripe[7867] = 24'h000000;
assign target_only_stripe[7868] = 24'h000000;
assign target_only_stripe[7869] = 24'h000000;
assign target_only_stripe[7870] = 24'h000000;
assign target_only_stripe[7871] = 24'h000000;
assign target_only_stripe[7872] = 24'h000000;
assign target_only_stripe[7873] = 24'h000000;
assign target_only_stripe[7874] = 24'h000000;
assign target_only_stripe[7875] = 24'h000000;
assign target_only_stripe[7876] = 24'h000000;
assign target_only_stripe[7877] = 24'h000000;
assign target_only_stripe[7878] = 24'h000000;
assign target_only_stripe[7879] = 24'h000000;
assign target_only_stripe[7880] = 24'h000000;
assign target_only_stripe[7881] = 24'h000000;
assign target_only_stripe[7882] = 24'h000000;
assign target_only_stripe[7883] = 24'h000000;
assign target_only_stripe[7884] = 24'h000000;
assign target_only_stripe[7885] = 24'h000000;
assign target_only_stripe[7886] = 24'h000000;
assign target_only_stripe[7887] = 24'h000000;
assign target_only_stripe[7888] = 24'h000000;
assign target_only_stripe[7889] = 24'h000000;
assign target_only_stripe[7890] = 24'h000000;
assign target_only_stripe[7891] = 24'h000000;
assign target_only_stripe[7892] = 24'h000000;
assign target_only_stripe[7893] = 24'h000000;
assign target_only_stripe[7894] = 24'h000000;
assign target_only_stripe[7895] = 24'h000000;
assign target_only_stripe[7896] = 24'h000000;
assign target_only_stripe[7897] = 24'h000000;
assign target_only_stripe[7898] = 24'h000000;
assign target_only_stripe[7899] = 24'h000000;
assign target_only_stripe[7900] = 24'h000000;
assign target_only_stripe[7901] = 24'h000000;
assign target_only_stripe[7902] = 24'h000000;
assign target_only_stripe[7903] = 24'h000000;
assign target_only_stripe[7904] = 24'h000000;
assign target_only_stripe[7905] = 24'h000000;
assign target_only_stripe[7906] = 24'h000000;
assign target_only_stripe[7907] = 24'h000000;
assign target_only_stripe[7908] = 24'h000000;
assign target_only_stripe[7909] = 24'h000000;
assign target_only_stripe[7910] = 24'h000000;
assign target_only_stripe[7911] = 24'h000000;
assign target_only_stripe[7912] = 24'h000000;
assign target_only_stripe[7913] = 24'h000000;
assign target_only_stripe[7914] = 24'h000000;
assign target_only_stripe[7915] = 24'h000000;
assign target_only_stripe[7916] = 24'h000000;
assign target_only_stripe[7917] = 24'h000000;
assign target_only_stripe[7918] = 24'h000000;
assign target_only_stripe[7919] = 24'h000000;
assign target_only_stripe[7920] = 24'h000000;
assign target_only_stripe[7921] = 24'h000000;
assign target_only_stripe[7922] = 24'h000000;
assign target_only_stripe[7923] = 24'h000000;
assign target_only_stripe[7924] = 24'h000000;
assign target_only_stripe[7925] = 24'h000000;
assign target_only_stripe[7926] = 24'h000000;
assign target_only_stripe[7927] = 24'h000000;
assign target_only_stripe[7928] = 24'hffffff;
assign target_only_stripe[7929] = 24'hffffff;
assign target_only_stripe[7930] = 24'hffffff;
assign target_only_stripe[7931] = 24'hffffff;
assign target_only_stripe[7932] = 24'hffffff;
assign target_only_stripe[7933] = 24'hffffff;
assign target_only_stripe[7934] = 24'hffffff;
assign target_only_stripe[7935] = 24'hffffff;
assign target_only_stripe[7936] = 24'hffffff;
assign target_only_stripe[7937] = 24'hffffff;
assign target_only_stripe[7938] = 24'hffffff;
assign target_only_stripe[7939] = 24'hffffff;
assign target_only_stripe[7940] = 24'hffffff;
assign target_only_stripe[7941] = 24'hffffff;
assign target_only_stripe[7942] = 24'hffffff;
assign target_only_stripe[7943] = 24'hffffff;
assign target_only_stripe[7944] = 24'hffffff;
assign target_only_stripe[7945] = 24'hffffff;
assign target_only_stripe[7946] = 24'hffffff;
assign target_only_stripe[7947] = 24'hffffff;
assign target_only_stripe[7948] = 24'hffffff;
assign target_only_stripe[7949] = 24'hffffff;
assign target_only_stripe[7950] = 24'hffffff;
assign target_only_stripe[7951] = 24'hffffff;
assign target_only_stripe[7952] = 24'hffffff;
assign target_only_stripe[7953] = 24'hffffff;
assign target_only_stripe[7954] = 24'hffffff;
assign target_only_stripe[7955] = 24'hffffff;
assign target_only_stripe[7956] = 24'hffffff;
assign target_only_stripe[7957] = 24'hffffff;
assign target_only_stripe[7958] = 24'hffffff;
assign target_only_stripe[7959] = 24'hffffff;
assign target_only_stripe[7960] = 24'hffffff;
assign target_only_stripe[7961] = 24'hffffff;
assign target_only_stripe[7962] = 24'hcccccc;
assign target_only_stripe[7963] = 24'h000000;
assign target_only_stripe[7964] = 24'h000000;
assign target_only_stripe[7965] = 24'h000000;
assign target_only_stripe[7966] = 24'h000000;
assign target_only_stripe[7967] = 24'h000000;
assign target_only_stripe[7968] = 24'h000000;
assign target_only_stripe[7969] = 24'h000000;
assign target_only_stripe[7970] = 24'h000000;
assign target_only_stripe[7971] = 24'h000000;
assign target_only_stripe[7972] = 24'h000000;
assign target_only_stripe[7973] = 24'h000000;
assign target_only_stripe[7974] = 24'h000000;
assign target_only_stripe[7975] = 24'h000000;
assign target_only_stripe[7976] = 24'h000000;
assign target_only_stripe[7977] = 24'h000000;
assign target_only_stripe[7978] = 24'h000000;
assign target_only_stripe[7979] = 24'h000000;
assign target_only_stripe[7980] = 24'h000000;
assign target_only_stripe[7981] = 24'h000000;
assign target_only_stripe[7982] = 24'h000000;
assign target_only_stripe[7983] = 24'h000000;
assign target_only_stripe[7984] = 24'h000000;
assign target_only_stripe[7985] = 24'h000000;
assign target_only_stripe[7986] = 24'h000000;
assign target_only_stripe[7987] = 24'h000000;
assign target_only_stripe[7988] = 24'h000000;
assign target_only_stripe[7989] = 24'h000000;
assign target_only_stripe[7990] = 24'h000000;
assign target_only_stripe[7991] = 24'h000000;
assign target_only_stripe[7992] = 24'h000000;
assign target_only_stripe[7993] = 24'h000000;
assign target_only_stripe[7994] = 24'h000000;
assign target_only_stripe[7995] = 24'hffffff;
assign target_only_stripe[7996] = 24'hffffff;
assign target_only_stripe[7997] = 24'hffffff;
assign target_only_stripe[7998] = 24'hffffff;
assign target_only_stripe[7999] = 24'hffffff;
assign target_only_stripe[8000] = 24'hffffff;
assign target_only_stripe[8001] = 24'hffffff;
assign target_only_stripe[8002] = 24'hffffff;
assign target_only_stripe[8003] = 24'hffffff;
assign target_only_stripe[8004] = 24'hffffff;
assign target_only_stripe[8005] = 24'hffffff;
assign target_only_stripe[8006] = 24'hffffff;
assign target_only_stripe[8007] = 24'hffffff;
assign target_only_stripe[8008] = 24'hffffff;
assign target_only_stripe[8009] = 24'hffffff;
assign target_only_stripe[8010] = 24'hffffff;
assign target_only_stripe[8011] = 24'hffffff;
assign target_only_stripe[8012] = 24'hffffff;
assign target_only_stripe[8013] = 24'hffffff;
assign target_only_stripe[8014] = 24'hffffff;
assign target_only_stripe[8015] = 24'hffffff;
assign target_only_stripe[8016] = 24'hffffff;
assign target_only_stripe[8017] = 24'hffffff;
assign target_only_stripe[8018] = 24'hffffff;
assign target_only_stripe[8019] = 24'hffffff;
assign target_only_stripe[8020] = 24'hffffff;
assign target_only_stripe[8021] = 24'hffffff;
assign target_only_stripe[8022] = 24'hffffff;
assign target_only_stripe[8023] = 24'hffffff;
assign target_only_stripe[8024] = 24'hffffff;
assign target_only_stripe[8025] = 24'hffffff;
assign target_only_stripe[8026] = 24'hffffff;
assign target_only_stripe[8027] = 24'hffffff;
assign target_only_stripe[8028] = 24'hffffff;
assign target_only_stripe[8029] = 24'hffffff;
assign target_only_stripe[8030] = 24'hffffff;
assign target_only_stripe[8031] = 24'h343434;
assign target_only_stripe[8032] = 24'h000000;
assign target_only_stripe[8033] = 24'h000000;
assign target_only_stripe[8034] = 24'h000000;
assign target_only_stripe[8035] = 24'h000000;
assign target_only_stripe[8036] = 24'h000000;
assign target_only_stripe[8037] = 24'h000000;
assign target_only_stripe[8038] = 24'h000000;
assign target_only_stripe[8039] = 24'h000000;
assign target_only_stripe[8040] = 24'h000000;
assign target_only_stripe[8041] = 24'h000000;
assign target_only_stripe[8042] = 24'h000000;
assign target_only_stripe[8043] = 24'h000000;
assign target_only_stripe[8044] = 24'h000000;
assign target_only_stripe[8045] = 24'h000000;
assign target_only_stripe[8046] = 24'h000000;
assign target_only_stripe[8047] = 24'h000000;
assign target_only_stripe[8048] = 24'h000000;
assign target_only_stripe[8049] = 24'h000000;
assign target_only_stripe[8050] = 24'h000000;
assign target_only_stripe[8051] = 24'h000000;
assign target_only_stripe[8052] = 24'h000000;
assign target_only_stripe[8053] = 24'h000000;
assign target_only_stripe[8054] = 24'h000000;
assign target_only_stripe[8055] = 24'h000000;
assign target_only_stripe[8056] = 24'h000000;
assign target_only_stripe[8057] = 24'h000000;
assign target_only_stripe[8058] = 24'h000000;
assign target_only_stripe[8059] = 24'h000000;
assign target_only_stripe[8060] = 24'h000000;
assign target_only_stripe[8061] = 24'h000000;
assign target_only_stripe[8062] = 24'h000000;
assign target_only_stripe[8063] = 24'h000000;
assign target_only_stripe[8064] = 24'h000000;
assign target_only_stripe[8065] = 24'h000000;
assign target_only_stripe[8066] = 24'h000000;
assign target_only_stripe[8067] = 24'h000000;
assign target_only_stripe[8068] = 24'h000000;
assign target_only_stripe[8069] = 24'h000000;
assign target_only_stripe[8070] = 24'h000000;
assign target_only_stripe[8071] = 24'h000000;
assign target_only_stripe[8072] = 24'h000000;
assign target_only_stripe[8073] = 24'h000000;
assign target_only_stripe[8074] = 24'h000000;
assign target_only_stripe[8075] = 24'h000000;
assign target_only_stripe[8076] = 24'h000000;
assign target_only_stripe[8077] = 24'h000000;
assign target_only_stripe[8078] = 24'h000000;
assign target_only_stripe[8079] = 24'h000000;
assign target_only_stripe[8080] = 24'h000000;
assign target_only_stripe[8081] = 24'h000000;
assign target_only_stripe[8082] = 24'h000000;
assign target_only_stripe[8083] = 24'h000000;
assign target_only_stripe[8084] = 24'h000000;
assign target_only_stripe[8085] = 24'h000000;
assign target_only_stripe[8086] = 24'h000000;
assign target_only_stripe[8087] = 24'h000000;
assign target_only_stripe[8088] = 24'h000000;
assign target_only_stripe[8089] = 24'h2d2d2d;
assign target_only_stripe[8090] = 24'hffffff;
assign target_only_stripe[8091] = 24'hffffff;
assign target_only_stripe[8092] = 24'hffffff;
assign target_only_stripe[8093] = 24'hffffff;
assign target_only_stripe[8094] = 24'hffffff;
assign target_only_stripe[8095] = 24'hffffff;
assign target_only_stripe[8096] = 24'hffffff;
assign target_only_stripe[8097] = 24'hffffff;
assign target_only_stripe[8098] = 24'hffffff;
assign target_only_stripe[8099] = 24'hffffff;
assign target_only_stripe[8100] = 24'hffffff;
assign target_only_stripe[8101] = 24'hffffff;
assign target_only_stripe[8102] = 24'hffffff;
assign target_only_stripe[8103] = 24'hffffff;
assign target_only_stripe[8104] = 24'hffffff;
assign target_only_stripe[8105] = 24'hffffff;
assign target_only_stripe[8106] = 24'hffffff;
assign target_only_stripe[8107] = 24'hffffff;
assign target_only_stripe[8108] = 24'hffffff;
assign target_only_stripe[8109] = 24'hffffff;
assign target_only_stripe[8110] = 24'hffffff;
assign target_only_stripe[8111] = 24'hffffff;
assign target_only_stripe[8112] = 24'hffffff;
assign target_only_stripe[8113] = 24'hffffff;
assign target_only_stripe[8114] = 24'hffffff;
assign target_only_stripe[8115] = 24'hffffff;
assign target_only_stripe[8116] = 24'hffffff;
assign target_only_stripe[8117] = 24'hffffff;
assign target_only_stripe[8118] = 24'hffffff;
assign target_only_stripe[8119] = 24'hffffff;
assign target_only_stripe[8120] = 24'hffffff;
assign target_only_stripe[8121] = 24'hffffff;
assign target_only_stripe[8122] = 24'hffffff;
assign target_only_stripe[8123] = 24'hffffff;
assign target_only_stripe[8124] = 24'hffffff;
assign target_only_stripe[8125] = 24'hffffff;
assign target_only_stripe[8126] = 24'h000000;
assign target_only_stripe[8127] = 24'h000000;
assign target_only_stripe[8128] = 24'h000000;
assign target_only_stripe[8129] = 24'h000000;
assign target_only_stripe[8130] = 24'h000000;
assign target_only_stripe[8131] = 24'h000000;
assign target_only_stripe[8132] = 24'h000000;
assign target_only_stripe[8133] = 24'h000000;
assign target_only_stripe[8134] = 24'h000000;
assign target_only_stripe[8135] = 24'h000000;
assign target_only_stripe[8136] = 24'h000000;
assign target_only_stripe[8137] = 24'h000000;
assign target_only_stripe[8138] = 24'h000000;
assign target_only_stripe[8139] = 24'h000000;
assign target_only_stripe[8140] = 24'h000000;
assign target_only_stripe[8141] = 24'h000000;
assign target_only_stripe[8142] = 24'h000000;
assign target_only_stripe[8143] = 24'h000000;
assign target_only_stripe[8144] = 24'h000000;
assign target_only_stripe[8145] = 24'h000000;
assign target_only_stripe[8146] = 24'h000000;
assign target_only_stripe[8147] = 24'h000000;
assign target_only_stripe[8148] = 24'h000000;
assign target_only_stripe[8149] = 24'h000000;
assign target_only_stripe[8150] = 24'h000000;
assign target_only_stripe[8151] = 24'h000000;
assign target_only_stripe[8152] = 24'h000000;
assign target_only_stripe[8153] = 24'h000000;
assign target_only_stripe[8154] = 24'h000000;
assign target_only_stripe[8155] = 24'h000000;
assign target_only_stripe[8156] = 24'h000000;
assign target_only_stripe[8157] = 24'h000000;
assign target_only_stripe[8158] = 24'he1e1e1;
assign target_only_stripe[8159] = 24'hffffff;
assign target_only_stripe[8160] = 24'hffffff;
assign target_only_stripe[8161] = 24'hffffff;
assign target_only_stripe[8162] = 24'hffffff;
assign target_only_stripe[8163] = 24'hffffff;
assign target_only_stripe[8164] = 24'hffffff;
assign target_only_stripe[8165] = 24'hffffff;
assign target_only_stripe[8166] = 24'hffffff;
assign target_only_stripe[8167] = 24'hffffff;
assign target_only_stripe[8168] = 24'hffffff;
assign target_only_stripe[8169] = 24'hffffff;
assign target_only_stripe[8170] = 24'hffffff;
assign target_only_stripe[8171] = 24'hffffff;
assign target_only_stripe[8172] = 24'hffffff;
assign target_only_stripe[8173] = 24'hffffff;
assign target_only_stripe[8174] = 24'hffffff;
assign target_only_stripe[8175] = 24'hffffff;
assign target_only_stripe[8176] = 24'hffffff;
assign target_only_stripe[8177] = 24'hffffff;
assign target_only_stripe[8178] = 24'hffffff;
assign target_only_stripe[8179] = 24'hffffff;
assign target_only_stripe[8180] = 24'hffffff;
assign target_only_stripe[8181] = 24'hffffff;
assign target_only_stripe[8182] = 24'hffffff;
assign target_only_stripe[8183] = 24'hffffff;
assign target_only_stripe[8184] = 24'hffffff;
assign target_only_stripe[8185] = 24'hffffff;
assign target_only_stripe[8186] = 24'hffffff;
assign target_only_stripe[8187] = 24'hffffff;
assign target_only_stripe[8188] = 24'hffffff;
assign target_only_stripe[8189] = 24'hffffff;
assign target_only_stripe[8190] = 24'hffffff;
assign target_only_stripe[8191] = 24'hffffff;
assign target_only_stripe[8192] = 24'he9e9e9;
assign target_only_stripe[8193] = 24'h000000;
assign target_only_stripe[8194] = 24'h000000;
assign target_only_stripe[8195] = 24'h000000;
assign target_only_stripe[8196] = 24'h000000;
assign target_only_stripe[8197] = 24'h000000;
assign target_only_stripe[8198] = 24'h000000;
assign target_only_stripe[8199] = 24'h000000;
assign target_only_stripe[8200] = 24'h000000;
assign target_only_stripe[8201] = 24'h000000;
assign target_only_stripe[8202] = 24'h000000;
assign target_only_stripe[8203] = 24'h000000;
assign target_only_stripe[8204] = 24'h000000;
assign target_only_stripe[8205] = 24'h000000;
assign target_only_stripe[8206] = 24'h000000;
assign target_only_stripe[8207] = 24'h000000;
assign target_only_stripe[8208] = 24'h000000;
assign target_only_stripe[8209] = 24'h000000;
assign target_only_stripe[8210] = 24'h000000;
assign target_only_stripe[8211] = 24'h000000;
assign target_only_stripe[8212] = 24'h000000;
assign target_only_stripe[8213] = 24'h000000;
assign target_only_stripe[8214] = 24'h000000;
assign target_only_stripe[8215] = 24'h000000;
assign target_only_stripe[8216] = 24'h000000;
assign target_only_stripe[8217] = 24'h000000;
assign target_only_stripe[8218] = 24'h000000;
assign target_only_stripe[8219] = 24'h000000;
assign target_only_stripe[8220] = 24'h000000;
assign target_only_stripe[8221] = 24'h000000;
assign target_only_stripe[8222] = 24'h000000;
assign target_only_stripe[8223] = 24'h000000;
assign target_only_stripe[8224] = 24'h000000;
assign target_only_stripe[8225] = 24'h010101;
assign target_only_stripe[8226] = 24'h000000;
assign target_only_stripe[8227] = 24'h000000;
assign target_only_stripe[8228] = 24'h000000;
assign target_only_stripe[8229] = 24'h000000;
assign target_only_stripe[8230] = 24'h000000;
assign target_only_stripe[8231] = 24'h000000;
assign target_only_stripe[8232] = 24'h000000;
assign target_only_stripe[8233] = 24'h000000;
assign target_only_stripe[8234] = 24'h000000;
assign target_only_stripe[8235] = 24'h000000;
assign target_only_stripe[8236] = 24'h000000;
assign target_only_stripe[8237] = 24'h000000;
assign target_only_stripe[8238] = 24'h000000;
assign target_only_stripe[8239] = 24'h000000;
assign target_only_stripe[8240] = 24'h000000;
assign target_only_stripe[8241] = 24'h000000;
assign target_only_stripe[8242] = 24'h000000;
assign target_only_stripe[8243] = 24'h000000;
assign target_only_stripe[8244] = 24'h000000;
assign target_only_stripe[8245] = 24'h000000;
assign target_only_stripe[8246] = 24'h000000;
assign target_only_stripe[8247] = 24'h000000;
assign target_only_stripe[8248] = 24'h000000;
assign target_only_stripe[8249] = 24'h000000;
assign target_only_stripe[8250] = 24'h000000;
assign target_only_stripe[8251] = 24'h000000;
assign target_only_stripe[8252] = 24'h000000;
assign target_only_stripe[8253] = 24'h000000;
assign target_only_stripe[8254] = 24'h000000;
assign target_only_stripe[8255] = 24'h000000;
assign target_only_stripe[8256] = 24'h000000;
assign target_only_stripe[8257] = 24'hffffff;
assign target_only_stripe[8258] = 24'hffffff;
assign target_only_stripe[8259] = 24'hffffff;
assign target_only_stripe[8260] = 24'hffffff;
assign target_only_stripe[8261] = 24'hffffff;
assign target_only_stripe[8262] = 24'hffffff;
assign target_only_stripe[8263] = 24'hffffff;
assign target_only_stripe[8264] = 24'hffffff;
assign target_only_stripe[8265] = 24'hffffff;
assign target_only_stripe[8266] = 24'hffffff;
assign target_only_stripe[8267] = 24'hffffff;
assign target_only_stripe[8268] = 24'hffffff;
assign target_only_stripe[8269] = 24'hffffff;
assign target_only_stripe[8270] = 24'hffffff;
assign target_only_stripe[8271] = 24'hffffff;
assign target_only_stripe[8272] = 24'hffffff;
assign target_only_stripe[8273] = 24'hffffff;
assign target_only_stripe[8274] = 24'hffffff;
assign target_only_stripe[8275] = 24'hffffff;
assign target_only_stripe[8276] = 24'hffffff;
assign target_only_stripe[8277] = 24'hffffff;
assign target_only_stripe[8278] = 24'hffffff;
assign target_only_stripe[8279] = 24'hffffff;
assign target_only_stripe[8280] = 24'hffffff;
assign target_only_stripe[8281] = 24'hffffff;
assign target_only_stripe[8282] = 24'hffffff;
assign target_only_stripe[8283] = 24'hffffff;
assign target_only_stripe[8284] = 24'hffffff;
assign target_only_stripe[8285] = 24'hffffff;
assign target_only_stripe[8286] = 24'hffffff;
assign target_only_stripe[8287] = 24'hffffff;
assign target_only_stripe[8288] = 24'hffffff;
assign target_only_stripe[8289] = 24'hffffff;
assign target_only_stripe[8290] = 24'hffffff;
assign target_only_stripe[8291] = 24'ha7a7a7;
assign target_only_stripe[8292] = 24'h000000;
assign target_only_stripe[8293] = 24'h000000;
assign target_only_stripe[8294] = 24'h000000;
assign target_only_stripe[8295] = 24'h000000;
assign target_only_stripe[8296] = 24'h000000;
assign target_only_stripe[8297] = 24'h000000;
assign target_only_stripe[8298] = 24'h000000;
assign target_only_stripe[8299] = 24'h000000;
assign target_only_stripe[8300] = 24'h000000;
assign target_only_stripe[8301] = 24'h000000;
assign target_only_stripe[8302] = 24'h000000;
assign target_only_stripe[8303] = 24'h000000;
assign target_only_stripe[8304] = 24'h000000;
assign target_only_stripe[8305] = 24'h000000;
assign target_only_stripe[8306] = 24'h000000;
assign target_only_stripe[8307] = 24'h000000;
assign target_only_stripe[8308] = 24'h000000;
assign target_only_stripe[8309] = 24'h000000;
assign target_only_stripe[8310] = 24'h000000;
assign target_only_stripe[8311] = 24'h000000;
assign target_only_stripe[8312] = 24'h000000;
assign target_only_stripe[8313] = 24'h000000;
assign target_only_stripe[8314] = 24'h000000;
assign target_only_stripe[8315] = 24'h000000;
assign target_only_stripe[8316] = 24'h000000;
assign target_only_stripe[8317] = 24'h000000;
assign target_only_stripe[8318] = 24'h000000;
assign target_only_stripe[8319] = 24'h000000;
assign target_only_stripe[8320] = 24'h000000;
assign target_only_stripe[8321] = 24'h000000;
assign target_only_stripe[8322] = 24'h000000;
assign target_only_stripe[8323] = 24'h000000;
assign target_only_stripe[8324] = 24'h3b3b3b;
assign target_only_stripe[8325] = 24'hffffff;
assign target_only_stripe[8326] = 24'hffffff;
assign target_only_stripe[8327] = 24'hffffff;
assign target_only_stripe[8328] = 24'hffffff;
assign target_only_stripe[8329] = 24'hffffff;
assign target_only_stripe[8330] = 24'hffffff;
assign target_only_stripe[8331] = 24'hffffff;
assign target_only_stripe[8332] = 24'hffffff;
assign target_only_stripe[8333] = 24'hffffff;
assign target_only_stripe[8334] = 24'hffffff;
assign target_only_stripe[8335] = 24'hffffff;
assign target_only_stripe[8336] = 24'hffffff;
assign target_only_stripe[8337] = 24'hffffff;
assign target_only_stripe[8338] = 24'hffffff;
assign target_only_stripe[8339] = 24'hffffff;
assign target_only_stripe[8340] = 24'hffffff;
assign target_only_stripe[8341] = 24'hffffff;
assign target_only_stripe[8342] = 24'hffffff;
assign target_only_stripe[8343] = 24'hffffff;
assign target_only_stripe[8344] = 24'hffffff;
assign target_only_stripe[8345] = 24'hffffff;
assign target_only_stripe[8346] = 24'hffffff;
assign target_only_stripe[8347] = 24'hffffff;
assign target_only_stripe[8348] = 24'hffffff;
assign target_only_stripe[8349] = 24'hffffff;
assign target_only_stripe[8350] = 24'hffffff;
assign target_only_stripe[8351] = 24'hffffff;
assign target_only_stripe[8352] = 24'hffffff;
assign target_only_stripe[8353] = 24'hffffff;
assign target_only_stripe[8354] = 24'hffffff;
assign target_only_stripe[8355] = 24'hffffff;
assign target_only_stripe[8356] = 24'hffffff;
assign target_only_stripe[8357] = 24'hffffff;
assign target_only_stripe[8358] = 24'hffffff;
assign target_only_stripe[8359] = 24'hffffff;
assign target_only_stripe[8360] = 24'h9a9a9a;
assign target_only_stripe[8361] = 24'h000000;
assign target_only_stripe[8362] = 24'h000000;
assign target_only_stripe[8363] = 24'h000000;
assign target_only_stripe[8364] = 24'h000000;
assign target_only_stripe[8365] = 24'h000000;
assign target_only_stripe[8366] = 24'h000000;
assign target_only_stripe[8367] = 24'h000000;
assign target_only_stripe[8368] = 24'h000000;
assign target_only_stripe[8369] = 24'h000000;
assign target_only_stripe[8370] = 24'h000000;
assign target_only_stripe[8371] = 24'h000000;
assign target_only_stripe[8372] = 24'h000000;
assign target_only_stripe[8373] = 24'h000000;
assign target_only_stripe[8374] = 24'h000000;
assign target_only_stripe[8375] = 24'h000000;
assign target_only_stripe[8376] = 24'h000000;
assign target_only_stripe[8377] = 24'h000000;
assign target_only_stripe[8378] = 24'h000000;
assign target_only_stripe[8379] = 24'h000000;
assign target_only_stripe[8380] = 24'h000000;
assign target_only_stripe[8381] = 24'h000000;
assign target_only_stripe[8382] = 24'h000000;
assign target_only_stripe[8383] = 24'h000000;
assign target_only_stripe[8384] = 24'h000000;
assign target_only_stripe[8385] = 24'h000000;
assign target_only_stripe[8386] = 24'h000000;
assign target_only_stripe[8387] = 24'h000000;
assign target_only_stripe[8388] = 24'h000000;
assign target_only_stripe[8389] = 24'h000000;
assign target_only_stripe[8390] = 24'h000000;
assign target_only_stripe[8391] = 24'h000000;
assign target_only_stripe[8392] = 24'h000000;
assign target_only_stripe[8393] = 24'h000000;
assign target_only_stripe[8394] = 24'h000000;
assign target_only_stripe[8395] = 24'h000000;
assign target_only_stripe[8396] = 24'h000000;
assign target_only_stripe[8397] = 24'h000000;
assign target_only_stripe[8398] = 24'h000000;
assign target_only_stripe[8399] = 24'h000000;
assign target_only_stripe[8400] = 24'h000000;
assign target_only_stripe[8401] = 24'h000000;
assign target_only_stripe[8402] = 24'h000000;
assign target_only_stripe[8403] = 24'h000000;
assign target_only_stripe[8404] = 24'h000000;
assign target_only_stripe[8405] = 24'h000000;
assign target_only_stripe[8406] = 24'h000000;
assign target_only_stripe[8407] = 24'h000000;
assign target_only_stripe[8408] = 24'h000000;
assign target_only_stripe[8409] = 24'h000000;
assign target_only_stripe[8410] = 24'h000000;
assign target_only_stripe[8411] = 24'h000000;
assign target_only_stripe[8412] = 24'h000000;
assign target_only_stripe[8413] = 24'h000000;
assign target_only_stripe[8414] = 24'h000000;
assign target_only_stripe[8415] = 24'h000000;
assign target_only_stripe[8416] = 24'h000000;
assign target_only_stripe[8417] = 24'h000000;
assign target_only_stripe[8418] = 24'h939393;
assign target_only_stripe[8419] = 24'hffffff;
assign target_only_stripe[8420] = 24'hffffff;
assign target_only_stripe[8421] = 24'hffffff;
assign target_only_stripe[8422] = 24'hffffff;
assign target_only_stripe[8423] = 24'hffffff;
assign target_only_stripe[8424] = 24'hffffff;
assign target_only_stripe[8425] = 24'hffffff;
assign target_only_stripe[8426] = 24'hffffff;
assign target_only_stripe[8427] = 24'hffffff;
assign target_only_stripe[8428] = 24'hffffff;
assign target_only_stripe[8429] = 24'hffffff;
assign target_only_stripe[8430] = 24'hffffff;
assign target_only_stripe[8431] = 24'hffffff;
assign target_only_stripe[8432] = 24'hffffff;
assign target_only_stripe[8433] = 24'hffffff;
assign target_only_stripe[8434] = 24'hffffff;
assign target_only_stripe[8435] = 24'hffffff;
assign target_only_stripe[8436] = 24'hffffff;
assign target_only_stripe[8437] = 24'hffffff;
assign target_only_stripe[8438] = 24'hffffff;
assign target_only_stripe[8439] = 24'hffffff;
assign target_only_stripe[8440] = 24'hffffff;
assign target_only_stripe[8441] = 24'hffffff;
assign target_only_stripe[8442] = 24'hffffff;
assign target_only_stripe[8443] = 24'hffffff;
assign target_only_stripe[8444] = 24'hffffff;
assign target_only_stripe[8445] = 24'hffffff;
assign target_only_stripe[8446] = 24'hffffff;
assign target_only_stripe[8447] = 24'hffffff;
assign target_only_stripe[8448] = 24'hffffff;
assign target_only_stripe[8449] = 24'hffffff;
assign target_only_stripe[8450] = 24'hffffff;
assign target_only_stripe[8451] = 24'hffffff;
assign target_only_stripe[8452] = 24'hffffff;
assign target_only_stripe[8453] = 24'hffffff;
assign target_only_stripe[8454] = 24'h454545;
assign target_only_stripe[8455] = 24'h000000;
assign target_only_stripe[8456] = 24'h000000;
assign target_only_stripe[8457] = 24'h000000;
assign target_only_stripe[8458] = 24'h000000;
assign target_only_stripe[8459] = 24'h000000;
assign target_only_stripe[8460] = 24'h000000;
assign target_only_stripe[8461] = 24'h000000;
assign target_only_stripe[8462] = 24'h000000;
assign target_only_stripe[8463] = 24'h000000;
assign target_only_stripe[8464] = 24'h000000;
assign target_only_stripe[8465] = 24'h000000;
assign target_only_stripe[8466] = 24'h000000;
assign target_only_stripe[8467] = 24'h000000;
assign target_only_stripe[8468] = 24'h000000;
assign target_only_stripe[8469] = 24'h000000;
assign target_only_stripe[8470] = 24'h000000;
assign target_only_stripe[8471] = 24'h000000;
assign target_only_stripe[8472] = 24'h000000;
assign target_only_stripe[8473] = 24'h000000;
assign target_only_stripe[8474] = 24'h000000;
assign target_only_stripe[8475] = 24'h000000;
assign target_only_stripe[8476] = 24'h000000;
assign target_only_stripe[8477] = 24'h000000;
assign target_only_stripe[8478] = 24'h000000;
assign target_only_stripe[8479] = 24'h000000;
assign target_only_stripe[8480] = 24'h000000;
assign target_only_stripe[8481] = 24'h000000;
assign target_only_stripe[8482] = 24'h000000;
assign target_only_stripe[8483] = 24'h000000;
assign target_only_stripe[8484] = 24'h000000;
assign target_only_stripe[8485] = 24'h000000;
assign target_only_stripe[8486] = 24'h000000;
assign target_only_stripe[8487] = 24'ha0a0a0;
assign target_only_stripe[8488] = 24'hffffff;
assign target_only_stripe[8489] = 24'hffffff;
assign target_only_stripe[8490] = 24'hffffff;
assign target_only_stripe[8491] = 24'hffffff;
assign target_only_stripe[8492] = 24'hffffff;
assign target_only_stripe[8493] = 24'hffffff;
assign target_only_stripe[8494] = 24'hffffff;
assign target_only_stripe[8495] = 24'hffffff;
assign target_only_stripe[8496] = 24'hffffff;
assign target_only_stripe[8497] = 24'hffffff;
assign target_only_stripe[8498] = 24'hffffff;
assign target_only_stripe[8499] = 24'hffffff;
assign target_only_stripe[8500] = 24'hffffff;
assign target_only_stripe[8501] = 24'hffffff;
assign target_only_stripe[8502] = 24'hffffff;
assign target_only_stripe[8503] = 24'hffffff;
assign target_only_stripe[8504] = 24'hffffff;
assign target_only_stripe[8505] = 24'hffffff;
assign target_only_stripe[8506] = 24'hffffff;
assign target_only_stripe[8507] = 24'hffffff;
assign target_only_stripe[8508] = 24'hffffff;
assign target_only_stripe[8509] = 24'hffffff;
assign target_only_stripe[8510] = 24'hffffff;
assign target_only_stripe[8511] = 24'hffffff;
assign target_only_stripe[8512] = 24'hffffff;
assign target_only_stripe[8513] = 24'hffffff;
assign target_only_stripe[8514] = 24'hffffff;
assign target_only_stripe[8515] = 24'hffffff;
assign target_only_stripe[8516] = 24'hffffff;
assign target_only_stripe[8517] = 24'hffffff;
assign target_only_stripe[8518] = 24'hffffff;
assign target_only_stripe[8519] = 24'hffffff;
assign target_only_stripe[8520] = 24'hffffff;
assign target_only_stripe[8521] = 24'hffffff;
assign target_only_stripe[8522] = 24'h000000;
assign target_only_stripe[8523] = 24'h000000;
assign target_only_stripe[8524] = 24'h000000;
assign target_only_stripe[8525] = 24'h000000;
assign target_only_stripe[8526] = 24'h000000;
assign target_only_stripe[8527] = 24'h000000;
assign target_only_stripe[8528] = 24'h000000;
assign target_only_stripe[8529] = 24'h000000;
assign target_only_stripe[8530] = 24'h000000;
assign target_only_stripe[8531] = 24'h000000;
assign target_only_stripe[8532] = 24'h000000;
assign target_only_stripe[8533] = 24'h000000;
assign target_only_stripe[8534] = 24'h000000;
assign target_only_stripe[8535] = 24'h000000;
assign target_only_stripe[8536] = 24'h000000;
assign target_only_stripe[8537] = 24'h000000;
assign target_only_stripe[8538] = 24'h000000;
assign target_only_stripe[8539] = 24'h000000;
assign target_only_stripe[8540] = 24'h000000;
assign target_only_stripe[8541] = 24'h000000;
assign target_only_stripe[8542] = 24'h000000;
assign target_only_stripe[8543] = 24'h000000;
assign target_only_stripe[8544] = 24'h000000;
assign target_only_stripe[8545] = 24'h000000;
assign target_only_stripe[8546] = 24'h000000;
assign target_only_stripe[8547] = 24'h000000;
assign target_only_stripe[8548] = 24'h000000;
assign target_only_stripe[8549] = 24'h000000;
assign target_only_stripe[8550] = 24'h000000;
assign target_only_stripe[8551] = 24'h000000;
assign target_only_stripe[8552] = 24'h000000;
assign target_only_stripe[8553] = 24'h000000;
assign target_only_stripe[8554] = 24'h010101;
assign target_only_stripe[8555] = 24'h000000;
assign target_only_stripe[8556] = 24'h000000;
assign target_only_stripe[8557] = 24'h000000;
assign target_only_stripe[8558] = 24'h000000;
assign target_only_stripe[8559] = 24'h000000;
assign target_only_stripe[8560] = 24'h000000;
assign target_only_stripe[8561] = 24'h000000;
assign target_only_stripe[8562] = 24'h000000;
assign target_only_stripe[8563] = 24'h000000;
assign target_only_stripe[8564] = 24'h000000;
assign target_only_stripe[8565] = 24'h000000;
assign target_only_stripe[8566] = 24'h000000;
assign target_only_stripe[8567] = 24'h000000;
assign target_only_stripe[8568] = 24'h000000;
assign target_only_stripe[8569] = 24'h000000;
assign target_only_stripe[8570] = 24'h000000;
assign target_only_stripe[8571] = 24'h000000;
assign target_only_stripe[8572] = 24'h000000;
assign target_only_stripe[8573] = 24'h000000;
assign target_only_stripe[8574] = 24'h000000;
assign target_only_stripe[8575] = 24'h000000;
assign target_only_stripe[8576] = 24'h000000;
assign target_only_stripe[8577] = 24'h000000;
assign target_only_stripe[8578] = 24'h000000;
assign target_only_stripe[8579] = 24'h000000;
assign target_only_stripe[8580] = 24'h000000;
assign target_only_stripe[8581] = 24'h000000;
assign target_only_stripe[8582] = 24'h000000;
assign target_only_stripe[8583] = 24'h000000;
assign target_only_stripe[8584] = 24'h000000;
assign target_only_stripe[8585] = 24'h000000;
assign target_only_stripe[8586] = 24'hffffff;
assign target_only_stripe[8587] = 24'hffffff;
assign target_only_stripe[8588] = 24'hffffff;
assign target_only_stripe[8589] = 24'hffffff;
assign target_only_stripe[8590] = 24'hffffff;
assign target_only_stripe[8591] = 24'hffffff;
assign target_only_stripe[8592] = 24'hffffff;
assign target_only_stripe[8593] = 24'hffffff;
assign target_only_stripe[8594] = 24'hffffff;
assign target_only_stripe[8595] = 24'hffffff;
assign target_only_stripe[8596] = 24'hffffff;
assign target_only_stripe[8597] = 24'hffffff;
assign target_only_stripe[8598] = 24'hffffff;
assign target_only_stripe[8599] = 24'hffffff;
assign target_only_stripe[8600] = 24'hffffff;
assign target_only_stripe[8601] = 24'hffffff;
assign target_only_stripe[8602] = 24'hffffff;
assign target_only_stripe[8603] = 24'hffffff;
assign target_only_stripe[8604] = 24'hffffff;
assign target_only_stripe[8605] = 24'hffffff;
assign target_only_stripe[8606] = 24'hffffff;
assign target_only_stripe[8607] = 24'hffffff;
assign target_only_stripe[8608] = 24'hffffff;
assign target_only_stripe[8609] = 24'hffffff;
assign target_only_stripe[8610] = 24'hffffff;
assign target_only_stripe[8611] = 24'hffffff;
assign target_only_stripe[8612] = 24'hffffff;
assign target_only_stripe[8613] = 24'hffffff;
assign target_only_stripe[8614] = 24'hffffff;
assign target_only_stripe[8615] = 24'hffffff;
assign target_only_stripe[8616] = 24'hffffff;
assign target_only_stripe[8617] = 24'hffffff;
assign target_only_stripe[8618] = 24'hffffff;
assign target_only_stripe[8619] = 24'hffffff;
assign target_only_stripe[8620] = 24'hc0c0c0;
assign target_only_stripe[8621] = 24'h010101;
assign target_only_stripe[8622] = 24'h000000;
assign target_only_stripe[8623] = 24'h000000;
assign target_only_stripe[8624] = 24'h000000;
assign target_only_stripe[8625] = 24'h000000;
assign target_only_stripe[8626] = 24'h000000;
assign target_only_stripe[8627] = 24'h000000;
assign target_only_stripe[8628] = 24'h000000;
assign target_only_stripe[8629] = 24'h000000;
assign target_only_stripe[8630] = 24'h000000;
assign target_only_stripe[8631] = 24'h000000;
assign target_only_stripe[8632] = 24'h000000;
assign target_only_stripe[8633] = 24'h000000;
assign target_only_stripe[8634] = 24'h000000;
assign target_only_stripe[8635] = 24'h000000;
assign target_only_stripe[8636] = 24'h000000;
assign target_only_stripe[8637] = 24'h000000;
assign target_only_stripe[8638] = 24'h000000;
assign target_only_stripe[8639] = 24'h000000;
assign target_only_stripe[8640] = 24'h000000;
assign target_only_stripe[8641] = 24'h000000;
assign target_only_stripe[8642] = 24'h000000;
assign target_only_stripe[8643] = 24'h000000;
assign target_only_stripe[8644] = 24'h000000;
assign target_only_stripe[8645] = 24'h000000;
assign target_only_stripe[8646] = 24'h000000;
assign target_only_stripe[8647] = 24'h000000;
assign target_only_stripe[8648] = 24'h000000;
assign target_only_stripe[8649] = 24'h000000;
assign target_only_stripe[8650] = 24'h000000;
assign target_only_stripe[8651] = 24'h000000;
assign target_only_stripe[8652] = 24'h000000;
assign target_only_stripe[8653] = 24'h121212;
assign target_only_stripe[8654] = 24'hffffff;
assign target_only_stripe[8655] = 24'hffffff;
assign target_only_stripe[8656] = 24'hffffff;
assign target_only_stripe[8657] = 24'hffffff;
assign target_only_stripe[8658] = 24'hffffff;
assign target_only_stripe[8659] = 24'hffffff;
assign target_only_stripe[8660] = 24'hffffff;
assign target_only_stripe[8661] = 24'hffffff;
assign target_only_stripe[8662] = 24'hffffff;
assign target_only_stripe[8663] = 24'hffffff;
assign target_only_stripe[8664] = 24'hffffff;
assign target_only_stripe[8665] = 24'hffffff;
assign target_only_stripe[8666] = 24'hffffff;
assign target_only_stripe[8667] = 24'hffffff;
assign target_only_stripe[8668] = 24'hffffff;
assign target_only_stripe[8669] = 24'hffffff;
assign target_only_stripe[8670] = 24'hffffff;
assign target_only_stripe[8671] = 24'hffffff;
assign target_only_stripe[8672] = 24'hffffff;
assign target_only_stripe[8673] = 24'hffffff;
assign target_only_stripe[8674] = 24'hffffff;
assign target_only_stripe[8675] = 24'hffffff;
assign target_only_stripe[8676] = 24'hffffff;
assign target_only_stripe[8677] = 24'hffffff;
assign target_only_stripe[8678] = 24'hffffff;
assign target_only_stripe[8679] = 24'hffffff;
assign target_only_stripe[8680] = 24'hffffff;
assign target_only_stripe[8681] = 24'hffffff;
assign target_only_stripe[8682] = 24'hffffff;
assign target_only_stripe[8683] = 24'hffffff;
assign target_only_stripe[8684] = 24'hffffff;
assign target_only_stripe[8685] = 24'hffffff;
assign target_only_stripe[8686] = 24'hffffff;
assign target_only_stripe[8687] = 24'hffffff;
assign target_only_stripe[8688] = 24'hffffff;
assign target_only_stripe[8689] = 24'hffffff;
assign target_only_stripe[8690] = 24'h343434;
assign target_only_stripe[8691] = 24'h000000;
assign target_only_stripe[8692] = 24'h000000;
assign target_only_stripe[8693] = 24'h000000;
assign target_only_stripe[8694] = 24'h000000;
assign target_only_stripe[8695] = 24'h000000;
assign target_only_stripe[8696] = 24'h000000;
assign target_only_stripe[8697] = 24'h000000;
assign target_only_stripe[8698] = 24'h000000;
assign target_only_stripe[8699] = 24'h000000;
assign target_only_stripe[8700] = 24'h000000;
assign target_only_stripe[8701] = 24'h000000;
assign target_only_stripe[8702] = 24'h000000;
assign target_only_stripe[8703] = 24'h000000;
assign target_only_stripe[8704] = 24'h000000;
assign target_only_stripe[8705] = 24'h000000;
assign target_only_stripe[8706] = 24'h000000;
assign target_only_stripe[8707] = 24'h000000;
assign target_only_stripe[8708] = 24'h000000;
assign target_only_stripe[8709] = 24'h000000;
assign target_only_stripe[8710] = 24'h000000;
assign target_only_stripe[8711] = 24'h000000;
assign target_only_stripe[8712] = 24'h000000;
assign target_only_stripe[8713] = 24'h000000;
assign target_only_stripe[8714] = 24'h000000;
assign target_only_stripe[8715] = 24'h000000;
assign target_only_stripe[8716] = 24'h000000;
assign target_only_stripe[8717] = 24'h000000;
assign target_only_stripe[8718] = 24'h000000;
assign target_only_stripe[8719] = 24'h000000;
assign target_only_stripe[8720] = 24'h000000;
assign target_only_stripe[8721] = 24'h000000;
assign target_only_stripe[8722] = 24'h000000;
assign target_only_stripe[8723] = 24'h000000;
assign target_only_stripe[8724] = 24'h000000;
assign target_only_stripe[8725] = 24'h000000;
assign target_only_stripe[8726] = 24'h000000;
assign target_only_stripe[8727] = 24'h000000;
assign target_only_stripe[8728] = 24'h000000;
assign target_only_stripe[8729] = 24'h000000;
assign target_only_stripe[8730] = 24'h000000;
assign target_only_stripe[8731] = 24'h000000;
assign target_only_stripe[8732] = 24'h000000;
assign target_only_stripe[8733] = 24'h000000;
assign target_only_stripe[8734] = 24'h000000;
assign target_only_stripe[8735] = 24'h000000;
assign target_only_stripe[8736] = 24'h000000;
assign target_only_stripe[8737] = 24'h000000;
assign target_only_stripe[8738] = 24'h000000;
assign target_only_stripe[8739] = 24'h000000;
assign target_only_stripe[8740] = 24'h000000;
assign target_only_stripe[8741] = 24'h000000;
assign target_only_stripe[8742] = 24'h000000;
assign target_only_stripe[8743] = 24'h000000;
assign target_only_stripe[8744] = 24'h000000;
assign target_only_stripe[8745] = 24'h000000;
assign target_only_stripe[8746] = 24'h2d2d2d;
assign target_only_stripe[8747] = 24'hffffff;
assign target_only_stripe[8748] = 24'hffffff;
assign target_only_stripe[8749] = 24'hffffff;
assign target_only_stripe[8750] = 24'hffffff;
assign target_only_stripe[8751] = 24'hffffff;
assign target_only_stripe[8752] = 24'hffffff;
assign target_only_stripe[8753] = 24'hffffff;
assign target_only_stripe[8754] = 24'hffffff;
assign target_only_stripe[8755] = 24'hffffff;
assign target_only_stripe[8756] = 24'hffffff;
assign target_only_stripe[8757] = 24'hffffff;
assign target_only_stripe[8758] = 24'hffffff;
assign target_only_stripe[8759] = 24'hffffff;
assign target_only_stripe[8760] = 24'hffffff;
assign target_only_stripe[8761] = 24'hffffff;
assign target_only_stripe[8762] = 24'hffffff;
assign target_only_stripe[8763] = 24'hffffff;
assign target_only_stripe[8764] = 24'hffffff;
assign target_only_stripe[8765] = 24'hffffff;
assign target_only_stripe[8766] = 24'hffffff;
assign target_only_stripe[8767] = 24'hffffff;
assign target_only_stripe[8768] = 24'hffffff;
assign target_only_stripe[8769] = 24'hffffff;
assign target_only_stripe[8770] = 24'hffffff;
assign target_only_stripe[8771] = 24'hffffff;
assign target_only_stripe[8772] = 24'hffffff;
assign target_only_stripe[8773] = 24'hffffff;
assign target_only_stripe[8774] = 24'hffffff;
assign target_only_stripe[8775] = 24'hffffff;
assign target_only_stripe[8776] = 24'hffffff;
assign target_only_stripe[8777] = 24'hffffff;
assign target_only_stripe[8778] = 24'hffffff;
assign target_only_stripe[8779] = 24'hffffff;
assign target_only_stripe[8780] = 24'hffffff;
assign target_only_stripe[8781] = 24'hffffff;
assign target_only_stripe[8782] = 24'hffffff;
assign target_only_stripe[8783] = 24'h171717;
assign target_only_stripe[8784] = 24'h000000;
assign target_only_stripe[8785] = 24'h000000;
assign target_only_stripe[8786] = 24'h000000;
assign target_only_stripe[8787] = 24'h000000;
assign target_only_stripe[8788] = 24'h000000;
assign target_only_stripe[8789] = 24'h000000;
assign target_only_stripe[8790] = 24'h000000;
assign target_only_stripe[8791] = 24'h000000;
assign target_only_stripe[8792] = 24'h000000;
assign target_only_stripe[8793] = 24'h000000;
assign target_only_stripe[8794] = 24'h000000;
assign target_only_stripe[8795] = 24'h000000;
assign target_only_stripe[8796] = 24'h000000;
assign target_only_stripe[8797] = 24'h000000;
assign target_only_stripe[8798] = 24'h000000;
assign target_only_stripe[8799] = 24'h000000;
assign target_only_stripe[8800] = 24'h000000;
assign target_only_stripe[8801] = 24'h000000;
assign target_only_stripe[8802] = 24'h000000;
assign target_only_stripe[8803] = 24'h000000;
assign target_only_stripe[8804] = 24'h000000;
assign target_only_stripe[8805] = 24'h000000;
assign target_only_stripe[8806] = 24'h000000;
assign target_only_stripe[8807] = 24'h000000;
assign target_only_stripe[8808] = 24'h000000;
assign target_only_stripe[8809] = 24'h000000;
assign target_only_stripe[8810] = 24'h000000;
assign target_only_stripe[8811] = 24'h000000;
assign target_only_stripe[8812] = 24'h000000;
assign target_only_stripe[8813] = 24'h000000;
assign target_only_stripe[8814] = 24'h000000;
assign target_only_stripe[8815] = 24'h010101;
assign target_only_stripe[8816] = 24'hbababa;
assign target_only_stripe[8817] = 24'hffffff;
assign target_only_stripe[8818] = 24'hffffff;
assign target_only_stripe[8819] = 24'hffffff;
assign target_only_stripe[8820] = 24'hffffff;
assign target_only_stripe[8821] = 24'hffffff;
assign target_only_stripe[8822] = 24'hffffff;
assign target_only_stripe[8823] = 24'hffffff;
assign target_only_stripe[8824] = 24'hffffff;
assign target_only_stripe[8825] = 24'hffffff;
assign target_only_stripe[8826] = 24'hffffff;
assign target_only_stripe[8827] = 24'hffffff;
assign target_only_stripe[8828] = 24'hffffff;
assign target_only_stripe[8829] = 24'hffffff;
assign target_only_stripe[8830] = 24'hffffff;
assign target_only_stripe[8831] = 24'hffffff;
assign target_only_stripe[8832] = 24'hffffff;
assign target_only_stripe[8833] = 24'hffffff;
assign target_only_stripe[8834] = 24'hffffff;
assign target_only_stripe[8835] = 24'hffffff;
assign target_only_stripe[8836] = 24'hffffff;
assign target_only_stripe[8837] = 24'hffffff;
assign target_only_stripe[8838] = 24'hffffff;
assign target_only_stripe[8839] = 24'hffffff;
assign target_only_stripe[8840] = 24'hffffff;
assign target_only_stripe[8841] = 24'hffffff;
assign target_only_stripe[8842] = 24'hffffff;
assign target_only_stripe[8843] = 24'hffffff;
assign target_only_stripe[8844] = 24'hffffff;
assign target_only_stripe[8845] = 24'hffffff;
assign target_only_stripe[8846] = 24'hffffff;
assign target_only_stripe[8847] = 24'hffffff;
assign target_only_stripe[8848] = 24'hffffff;
assign target_only_stripe[8849] = 24'hffffff;
assign target_only_stripe[8850] = 24'hffffff;
assign target_only_stripe[8851] = 24'h000000;
assign target_only_stripe[8852] = 24'h000000;
assign target_only_stripe[8853] = 24'h000000;
assign target_only_stripe[8854] = 24'h000000;
assign target_only_stripe[8855] = 24'h000000;
assign target_only_stripe[8856] = 24'h000000;
assign target_only_stripe[8857] = 24'h000000;
assign target_only_stripe[8858] = 24'h000000;
assign target_only_stripe[8859] = 24'h000000;
assign target_only_stripe[8860] = 24'h000000;
assign target_only_stripe[8861] = 24'h000000;
assign target_only_stripe[8862] = 24'h000000;
assign target_only_stripe[8863] = 24'h000000;
assign target_only_stripe[8864] = 24'h000000;
assign target_only_stripe[8865] = 24'h000000;
assign target_only_stripe[8866] = 24'h000000;
assign target_only_stripe[8867] = 24'h000000;
assign target_only_stripe[8868] = 24'h000000;
assign target_only_stripe[8869] = 24'h000000;
assign target_only_stripe[8870] = 24'h000000;
assign target_only_stripe[8871] = 24'h000000;
assign target_only_stripe[8872] = 24'h000000;
assign target_only_stripe[8873] = 24'h000000;
assign target_only_stripe[8874] = 24'h000000;
assign target_only_stripe[8875] = 24'h000000;
assign target_only_stripe[8876] = 24'h000000;
assign target_only_stripe[8877] = 24'h000000;
assign target_only_stripe[8878] = 24'h000000;
assign target_only_stripe[8879] = 24'h000000;
assign target_only_stripe[8880] = 24'h000000;
assign target_only_stripe[8881] = 24'h000000;
assign target_only_stripe[8882] = 24'h000000;
assign target_only_stripe[8883] = 24'h070707;
assign target_only_stripe[8884] = 24'h000000;
assign target_only_stripe[8885] = 24'h000000;
assign target_only_stripe[8886] = 24'h000000;
assign target_only_stripe[8887] = 24'h000000;
assign target_only_stripe[8888] = 24'h000000;
assign target_only_stripe[8889] = 24'h000000;
assign target_only_stripe[8890] = 24'h000000;
assign target_only_stripe[8891] = 24'h000000;
assign target_only_stripe[8892] = 24'h000000;
assign target_only_stripe[8893] = 24'h000000;
assign target_only_stripe[8894] = 24'h000000;
assign target_only_stripe[8895] = 24'h000000;
assign target_only_stripe[8896] = 24'h000000;
assign target_only_stripe[8897] = 24'h000000;
assign target_only_stripe[8898] = 24'h000000;
assign target_only_stripe[8899] = 24'h000000;
assign target_only_stripe[8900] = 24'h000000;
assign target_only_stripe[8901] = 24'h000000;
assign target_only_stripe[8902] = 24'h000000;
assign target_only_stripe[8903] = 24'h000000;
assign target_only_stripe[8904] = 24'h000000;
assign target_only_stripe[8905] = 24'h000000;
assign target_only_stripe[8906] = 24'h000000;
assign target_only_stripe[8907] = 24'h000000;
assign target_only_stripe[8908] = 24'h000000;
assign target_only_stripe[8909] = 24'h000000;
assign target_only_stripe[8910] = 24'h000000;
assign target_only_stripe[8911] = 24'h000000;
assign target_only_stripe[8912] = 24'h000000;
assign target_only_stripe[8913] = 24'h000000;
assign target_only_stripe[8914] = 24'h000000;
assign target_only_stripe[8915] = 24'h999999;
assign target_only_stripe[8916] = 24'hd6c9c4;
assign target_only_stripe[8917] = 24'hffffff;
assign target_only_stripe[8918] = 24'hffffff;
assign target_only_stripe[8919] = 24'hffffff;
assign target_only_stripe[8920] = 24'hffffff;
assign target_only_stripe[8921] = 24'hffffff;
assign target_only_stripe[8922] = 24'hffffff;
assign target_only_stripe[8923] = 24'hffffff;
assign target_only_stripe[8924] = 24'hffffff;
assign target_only_stripe[8925] = 24'hffffff;
assign target_only_stripe[8926] = 24'hffffff;
assign target_only_stripe[8927] = 24'hffffff;
assign target_only_stripe[8928] = 24'hffffff;
assign target_only_stripe[8929] = 24'hffffff;
assign target_only_stripe[8930] = 24'hffffff;
assign target_only_stripe[8931] = 24'hffffff;
assign target_only_stripe[8932] = 24'hffffff;
assign target_only_stripe[8933] = 24'hffffff;
assign target_only_stripe[8934] = 24'hffffff;
assign target_only_stripe[8935] = 24'hffffff;
assign target_only_stripe[8936] = 24'hffffff;
assign target_only_stripe[8937] = 24'hffffff;
assign target_only_stripe[8938] = 24'hffffff;
assign target_only_stripe[8939] = 24'hffffff;
assign target_only_stripe[8940] = 24'hffffff;
assign target_only_stripe[8941] = 24'hffffff;
assign target_only_stripe[8942] = 24'hffffff;
assign target_only_stripe[8943] = 24'hffffff;
assign target_only_stripe[8944] = 24'hffffff;
assign target_only_stripe[8945] = 24'hffffff;
assign target_only_stripe[8946] = 24'hffffff;
assign target_only_stripe[8947] = 24'hffffff;
assign target_only_stripe[8948] = 24'hffffff;
assign target_only_stripe[8949] = 24'hd7d7d7;
assign target_only_stripe[8950] = 24'h141414;
assign target_only_stripe[8951] = 24'h000000;
assign target_only_stripe[8952] = 24'h000000;
assign target_only_stripe[8953] = 24'h000000;
assign target_only_stripe[8954] = 24'h000000;
assign target_only_stripe[8955] = 24'h000000;
assign target_only_stripe[8956] = 24'h000000;
assign target_only_stripe[8957] = 24'h000000;
assign target_only_stripe[8958] = 24'h000000;
assign target_only_stripe[8959] = 24'h000000;
assign target_only_stripe[8960] = 24'h000000;
assign target_only_stripe[8961] = 24'h000000;
assign target_only_stripe[8962] = 24'h000000;
assign target_only_stripe[8963] = 24'h000000;
assign target_only_stripe[8964] = 24'h000000;
assign target_only_stripe[8965] = 24'h000000;
assign target_only_stripe[8966] = 24'h000000;
assign target_only_stripe[8967] = 24'h000000;
assign target_only_stripe[8968] = 24'h000000;
assign target_only_stripe[8969] = 24'h000000;
assign target_only_stripe[8970] = 24'h000000;
assign target_only_stripe[8971] = 24'h000000;
assign target_only_stripe[8972] = 24'h000000;
assign target_only_stripe[8973] = 24'h000000;
assign target_only_stripe[8974] = 24'h000000;
assign target_only_stripe[8975] = 24'h000000;
assign target_only_stripe[8976] = 24'h000000;
assign target_only_stripe[8977] = 24'h000000;
assign target_only_stripe[8978] = 24'h000000;
assign target_only_stripe[8979] = 24'h000000;
assign target_only_stripe[8980] = 24'h000000;
assign target_only_stripe[8981] = 24'h000000;
assign target_only_stripe[8982] = 24'h000000;
assign target_only_stripe[8983] = 24'ha3a3a3;
assign target_only_stripe[8984] = 24'hffffff;
assign target_only_stripe[8985] = 24'hffffff;
assign target_only_stripe[8986] = 24'hffffff;
assign target_only_stripe[8987] = 24'hffffff;
assign target_only_stripe[8988] = 24'hffffff;
assign target_only_stripe[8989] = 24'hffffff;
assign target_only_stripe[8990] = 24'hffffff;
assign target_only_stripe[8991] = 24'hffffff;
assign target_only_stripe[8992] = 24'hffffff;
assign target_only_stripe[8993] = 24'hffffff;
assign target_only_stripe[8994] = 24'hffffff;
assign target_only_stripe[8995] = 24'hffffff;
assign target_only_stripe[8996] = 24'hffffff;
assign target_only_stripe[8997] = 24'hffffff;
assign target_only_stripe[8998] = 24'hffffff;
assign target_only_stripe[8999] = 24'hffffff;
assign target_only_stripe[9000] = 24'hffffff;
assign target_only_stripe[9001] = 24'hffffff;
assign target_only_stripe[9002] = 24'hffffff;
assign target_only_stripe[9003] = 24'hffffff;
assign target_only_stripe[9004] = 24'hffffff;
assign target_only_stripe[9005] = 24'hffffff;
assign target_only_stripe[9006] = 24'hffffff;
assign target_only_stripe[9007] = 24'hffffff;
assign target_only_stripe[9008] = 24'hffffff;
assign target_only_stripe[9009] = 24'hffffff;
assign target_only_stripe[9010] = 24'hffffff;
assign target_only_stripe[9011] = 24'hffffff;
assign target_only_stripe[9012] = 24'hffffff;
assign target_only_stripe[9013] = 24'hffffff;
assign target_only_stripe[9014] = 24'hffffff;
assign target_only_stripe[9015] = 24'hffffff;
assign target_only_stripe[9016] = 24'hffffff;
assign target_only_stripe[9017] = 24'hffffff;
assign target_only_stripe[9018] = 24'hffffff;
assign target_only_stripe[9019] = 24'h9b9b9b;
assign target_only_stripe[9020] = 24'h010101;
assign target_only_stripe[9021] = 24'h000000;
assign target_only_stripe[9022] = 24'h000000;
assign target_only_stripe[9023] = 24'h000000;
assign target_only_stripe[9024] = 24'h000000;
assign target_only_stripe[9025] = 24'h000000;
assign target_only_stripe[9026] = 24'h000000;
assign target_only_stripe[9027] = 24'h000000;
assign target_only_stripe[9028] = 24'h000000;
assign target_only_stripe[9029] = 24'h000000;
assign target_only_stripe[9030] = 24'h000000;
assign target_only_stripe[9031] = 24'h000000;
assign target_only_stripe[9032] = 24'h000000;
assign target_only_stripe[9033] = 24'h000000;
assign target_only_stripe[9034] = 24'h000000;
assign target_only_stripe[9035] = 24'h000000;
assign target_only_stripe[9036] = 24'h000000;
assign target_only_stripe[9037] = 24'h000000;
assign target_only_stripe[9038] = 24'h000000;
assign target_only_stripe[9039] = 24'h000000;
assign target_only_stripe[9040] = 24'h000000;
assign target_only_stripe[9041] = 24'h000000;
assign target_only_stripe[9042] = 24'h000000;
assign target_only_stripe[9043] = 24'h000000;
assign target_only_stripe[9044] = 24'h000000;
assign target_only_stripe[9045] = 24'h000000;
assign target_only_stripe[9046] = 24'h000000;
assign target_only_stripe[9047] = 24'h000000;
assign target_only_stripe[9048] = 24'h000000;
assign target_only_stripe[9049] = 24'h000000;
assign target_only_stripe[9050] = 24'h000000;
assign target_only_stripe[9051] = 24'h000000;
assign target_only_stripe[9052] = 24'h000000;
assign target_only_stripe[9053] = 24'h000000;
assign target_only_stripe[9054] = 24'h000000;
assign target_only_stripe[9055] = 24'h000000;
assign target_only_stripe[9056] = 24'h000000;
assign target_only_stripe[9057] = 24'h000000;
assign target_only_stripe[9058] = 24'h000000;
assign target_only_stripe[9059] = 24'h000000;
assign target_only_stripe[9060] = 24'h000000;
assign target_only_stripe[9061] = 24'h000000;
assign target_only_stripe[9062] = 24'h000000;
assign target_only_stripe[9063] = 24'h000000;
assign target_only_stripe[9064] = 24'h000000;
assign target_only_stripe[9065] = 24'h000000;
assign target_only_stripe[9066] = 24'h000000;
assign target_only_stripe[9067] = 24'h000000;
assign target_only_stripe[9068] = 24'h000000;
assign target_only_stripe[9069] = 24'h000000;
assign target_only_stripe[9070] = 24'h000000;
assign target_only_stripe[9071] = 24'h000000;
assign target_only_stripe[9072] = 24'h000000;
assign target_only_stripe[9073] = 24'h000000;
assign target_only_stripe[9074] = 24'h010101;
assign target_only_stripe[9075] = 24'h949494;
assign target_only_stripe[9076] = 24'hffffff;
assign target_only_stripe[9077] = 24'hffffff;
assign target_only_stripe[9078] = 24'hffffff;
assign target_only_stripe[9079] = 24'hffffff;
assign target_only_stripe[9080] = 24'hffffff;
assign target_only_stripe[9081] = 24'hffffff;
assign target_only_stripe[9082] = 24'hffffff;
assign target_only_stripe[9083] = 24'hffffff;
assign target_only_stripe[9084] = 24'hffffff;
assign target_only_stripe[9085] = 24'hffffff;
assign target_only_stripe[9086] = 24'hffffff;
assign target_only_stripe[9087] = 24'hffffff;
assign target_only_stripe[9088] = 24'hffffff;
assign target_only_stripe[9089] = 24'hffffff;
assign target_only_stripe[9090] = 24'hffffff;
assign target_only_stripe[9091] = 24'hffffff;
assign target_only_stripe[9092] = 24'hffffff;
assign target_only_stripe[9093] = 24'hffffff;
assign target_only_stripe[9094] = 24'hffffff;
assign target_only_stripe[9095] = 24'hffffff;
assign target_only_stripe[9096] = 24'hffffff;
assign target_only_stripe[9097] = 24'hffffff;
assign target_only_stripe[9098] = 24'hffffff;
assign target_only_stripe[9099] = 24'hffffff;
assign target_only_stripe[9100] = 24'hffffff;
assign target_only_stripe[9101] = 24'hffffff;
assign target_only_stripe[9102] = 24'hffffff;
assign target_only_stripe[9103] = 24'hffffff;
assign target_only_stripe[9104] = 24'hffffff;
assign target_only_stripe[9105] = 24'hffffff;
assign target_only_stripe[9106] = 24'hffffff;
assign target_only_stripe[9107] = 24'hffffff;
assign target_only_stripe[9108] = 24'hffffff;
assign target_only_stripe[9109] = 24'hffffff;
assign target_only_stripe[9110] = 24'hffffff;
assign target_only_stripe[9111] = 24'haaaaaa;
assign target_only_stripe[9112] = 24'h000000;
assign target_only_stripe[9113] = 24'h000000;
assign target_only_stripe[9114] = 24'h000000;
assign target_only_stripe[9115] = 24'h000000;
assign target_only_stripe[9116] = 24'h000000;
assign target_only_stripe[9117] = 24'h000000;
assign target_only_stripe[9118] = 24'h000000;
assign target_only_stripe[9119] = 24'h000000;
assign target_only_stripe[9120] = 24'h000000;
assign target_only_stripe[9121] = 24'h000000;
assign target_only_stripe[9122] = 24'h000000;
assign target_only_stripe[9123] = 24'h000000;
assign target_only_stripe[9124] = 24'h000000;
assign target_only_stripe[9125] = 24'h000000;
assign target_only_stripe[9126] = 24'h000000;
assign target_only_stripe[9127] = 24'h000000;
assign target_only_stripe[9128] = 24'h000000;
assign target_only_stripe[9129] = 24'h000000;
assign target_only_stripe[9130] = 24'h000000;
assign target_only_stripe[9131] = 24'h000000;
assign target_only_stripe[9132] = 24'h000000;
assign target_only_stripe[9133] = 24'h000000;
assign target_only_stripe[9134] = 24'h000000;
assign target_only_stripe[9135] = 24'h000000;
assign target_only_stripe[9136] = 24'h000000;
assign target_only_stripe[9137] = 24'h000000;
assign target_only_stripe[9138] = 24'h000000;
assign target_only_stripe[9139] = 24'h000000;
assign target_only_stripe[9140] = 24'h000000;
assign target_only_stripe[9141] = 24'h000000;
assign target_only_stripe[9142] = 24'h000000;
assign target_only_stripe[9143] = 24'h000000;
assign target_only_stripe[9144] = 24'h0e0e0e;
assign target_only_stripe[9145] = 24'hd2d2d2;
assign target_only_stripe[9146] = 24'hffffff;
assign target_only_stripe[9147] = 24'hffffff;
assign target_only_stripe[9148] = 24'hffffff;
assign target_only_stripe[9149] = 24'hffffff;
assign target_only_stripe[9150] = 24'hffffff;
assign target_only_stripe[9151] = 24'hffffff;
assign target_only_stripe[9152] = 24'hffffff;
assign target_only_stripe[9153] = 24'hffffff;
assign target_only_stripe[9154] = 24'hffffff;
assign target_only_stripe[9155] = 24'hffffff;
assign target_only_stripe[9156] = 24'hffffff;
assign target_only_stripe[9157] = 24'hffffff;
assign target_only_stripe[9158] = 24'hffffff;
assign target_only_stripe[9159] = 24'hffffff;
assign target_only_stripe[9160] = 24'hffffff;
assign target_only_stripe[9161] = 24'hffffff;
assign target_only_stripe[9162] = 24'hffffff;
assign target_only_stripe[9163] = 24'hffffff;
assign target_only_stripe[9164] = 24'hffffff;
assign target_only_stripe[9165] = 24'hffffff;
assign target_only_stripe[9166] = 24'hffffff;
assign target_only_stripe[9167] = 24'hffffff;
assign target_only_stripe[9168] = 24'hffffff;
assign target_only_stripe[9169] = 24'hffffff;
assign target_only_stripe[9170] = 24'hffffff;
assign target_only_stripe[9171] = 24'hffffff;
assign target_only_stripe[9172] = 24'hffffff;
assign target_only_stripe[9173] = 24'hffffff;
assign target_only_stripe[9174] = 24'hffffff;
assign target_only_stripe[9175] = 24'hffffff;
assign target_only_stripe[9176] = 24'hffffff;
assign target_only_stripe[9177] = 24'hffffff;
assign target_only_stripe[9178] = 24'hffffff;
assign target_only_stripe[9179] = 24'hbdbdbd;
assign target_only_stripe[9180] = 24'h000000;
assign target_only_stripe[9181] = 24'h000000;
assign target_only_stripe[9182] = 24'h000000;
assign target_only_stripe[9183] = 24'h000000;
assign target_only_stripe[9184] = 24'h000000;
assign target_only_stripe[9185] = 24'h000000;
assign target_only_stripe[9186] = 24'h000000;
assign target_only_stripe[9187] = 24'h000000;
assign target_only_stripe[9188] = 24'h000000;
assign target_only_stripe[9189] = 24'h000000;
assign target_only_stripe[9190] = 24'h000000;
assign target_only_stripe[9191] = 24'h000000;
assign target_only_stripe[9192] = 24'h000000;
assign target_only_stripe[9193] = 24'h000000;
assign target_only_stripe[9194] = 24'h000000;
assign target_only_stripe[9195] = 24'h000000;
assign target_only_stripe[9196] = 24'h000000;
assign target_only_stripe[9197] = 24'h000000;
assign target_only_stripe[9198] = 24'h000000;
assign target_only_stripe[9199] = 24'h000000;
assign target_only_stripe[9200] = 24'h000000;
assign target_only_stripe[9201] = 24'h000000;
assign target_only_stripe[9202] = 24'h000000;
assign target_only_stripe[9203] = 24'h000000;
assign target_only_stripe[9204] = 24'h000000;
assign target_only_stripe[9205] = 24'h000000;
assign target_only_stripe[9206] = 24'h000000;
assign target_only_stripe[9207] = 24'h000000;
assign target_only_stripe[9208] = 24'h000000;
assign target_only_stripe[9209] = 24'h000000;
assign target_only_stripe[9210] = 24'h000000;
assign target_only_stripe[9211] = 24'h040404;
