localparam NUM_PIXELS_TARGET7 = 400;
logic [23:0] target7 [0:399];
assign target7[0] = 24'h000000;
assign target7[1] = 24'hffffff;
assign target7[2] = 24'h000000;
assign target7[3] = 24'hffffff;
assign target7[4] = 24'h000000;
assign target7[5] = 24'hffffff;
assign target7[6] = 24'h000000;
assign target7[7] = 24'hffffff;
assign target7[8] = 24'hff0000;
assign target7[9] = 24'hff0000;
assign target7[10] = 24'hffffff;
assign target7[11] = 24'hffffff;
assign target7[12] = 24'h00ff00;
assign target7[13] = 24'h00ff00;
assign target7[14] = 24'hffffff;
assign target7[15] = 24'hffffff;
assign target7[16] = 24'h0000ff;
assign target7[17] = 24'h0000ff;
assign target7[18] = 24'hffffff;
assign target7[19] = 24'hffffff;
assign target7[20] = 24'h00ffff;
assign target7[21] = 24'h00ffff;
assign target7[22] = 24'hffffff;
assign target7[23] = 24'hffffff;
assign target7[24] = 24'hff00ff;
assign target7[25] = 24'hff00ff;
assign target7[26] = 24'hffffff;
assign target7[27] = 24'hffffff;
assign target7[28] = 24'hffff00;
assign target7[29] = 24'hffff00;
assign target7[30] = 24'hffffff;
assign target7[31] = 24'hffffff;
assign target7[32] = 24'h000000;
assign target7[33] = 24'h000000;
assign target7[34] = 24'h000000;
assign target7[35] = 24'h000000;
assign target7[36] = 24'h000000;
assign target7[37] = 24'h000000;
assign target7[38] = 24'h000000;
assign target7[39] = 24'h000000;
assign target7[40] = 24'h8f8f8f;
assign target7[41] = 24'h8f8f8f;
assign target7[42] = 24'h8f8f8f;
assign target7[43] = 24'h8f8f8f;
assign target7[44] = 24'hffffff;
assign target7[45] = 24'hffffff;
assign target7[46] = 24'hffffff;
assign target7[47] = 24'hffffff;
assign target7[48] = 24'h8f8f8f;
assign target7[49] = 24'h8f8f8f;
assign target7[50] = 24'h8f8f8f;
assign target7[51] = 24'h8f8f8f;
assign target7[52] = 24'hffffff;
assign target7[53] = 24'hffffff;
assign target7[54] = 24'hffffff;
assign target7[55] = 24'hffffff;
assign target7[56] = 24'h000000;
assign target7[57] = 24'h000000;
assign target7[58] = 24'h000000;
assign target7[59] = 24'hffffff;
assign target7[60] = 24'hffffff;
assign target7[61] = 24'hffffff;
assign target7[62] = 24'hffffff;
assign target7[63] = 24'hffffff;
assign target7[64] = 24'hffffff;
assign target7[65] = 24'hffffff;
assign target7[66] = 24'hffffff;
assign target7[67] = 24'hffffff;
assign target7[68] = 24'hffffff;
assign target7[69] = 24'hffffff;
assign target7[70] = 24'hffffff;
assign target7[71] = 24'hffffff;
assign target7[72] = 24'hffffff;
assign target7[73] = 24'hffffff;
assign target7[74] = 24'hffffff;
assign target7[75] = 24'hffffff;
assign target7[76] = 24'hffffff;
assign target7[77] = 24'hffffff;
assign target7[78] = 24'hffffff;
assign target7[79] = 24'hffffff;
assign target7[80] = 24'h000000;
assign target7[81] = 24'h000000;
assign target7[82] = 24'h000000;
assign target7[83] = 24'h000000;
assign target7[84] = 24'h000000;
assign target7[85] = 24'h000000;
assign target7[86] = 24'h000000;
assign target7[87] = 24'h000000;
assign target7[88] = 24'h000000;
assign target7[89] = 24'h000000;
assign target7[90] = 24'h000000;
assign target7[91] = 24'h000000;
assign target7[92] = 24'h000000;
assign target7[93] = 24'h000000;
assign target7[94] = 24'h000000;
assign target7[95] = 24'h000000;
assign target7[96] = 24'h000000;
assign target7[97] = 24'h000000;
assign target7[98] = 24'h000000;
assign target7[99] = 24'h000000;
assign target7[100] = 24'hff0000;
assign target7[101] = 24'hff0000;
assign target7[102] = 24'hff0000;
assign target7[103] = 24'hff0000;
assign target7[104] = 24'hff0000;
assign target7[105] = 24'hff0000;
assign target7[106] = 24'hff0000;
assign target7[107] = 24'hff0000;
assign target7[108] = 24'hff0000;
assign target7[109] = 24'hff0000;
assign target7[110] = 24'hff0000;
assign target7[111] = 24'hff0000;
assign target7[112] = 24'hff0000;
assign target7[113] = 24'hff0000;
assign target7[114] = 24'hff0000;
assign target7[115] = 24'hff0000;
assign target7[116] = 24'hff0000;
assign target7[117] = 24'hff0000;
assign target7[118] = 24'hff0000;
assign target7[119] = 24'hff0000;
assign target7[120] = 24'h00ff00;
assign target7[121] = 24'h00ff00;
assign target7[122] = 24'h00ff00;
assign target7[123] = 24'h00ff00;
assign target7[124] = 24'h00ff00;
assign target7[125] = 24'h00ff00;
assign target7[126] = 24'h00ff00;
assign target7[127] = 24'h00ff00;
assign target7[128] = 24'h00ff00;
assign target7[129] = 24'h00ff00;
assign target7[130] = 24'h00ff00;
assign target7[131] = 24'h00ff00;
assign target7[132] = 24'h00ff00;
assign target7[133] = 24'h00ff00;
assign target7[134] = 24'h00ff00;
assign target7[135] = 24'h00ff00;
assign target7[136] = 24'h00ff00;
assign target7[137] = 24'h00ff00;
assign target7[138] = 24'h00ff00;
assign target7[139] = 24'h00ff00;
assign target7[140] = 24'h0000ff;
assign target7[141] = 24'h0000ff;
assign target7[142] = 24'h0000ff;
assign target7[143] = 24'h0000ff;
assign target7[144] = 24'h0000ff;
assign target7[145] = 24'h0000ff;
assign target7[146] = 24'h0000ff;
assign target7[147] = 24'h0000ff;
assign target7[148] = 24'h0000ff;
assign target7[149] = 24'h0000ff;
assign target7[150] = 24'h0000ff;
assign target7[151] = 24'h0000ff;
assign target7[152] = 24'h0000ff;
assign target7[153] = 24'h0000ff;
assign target7[154] = 24'h0000ff;
assign target7[155] = 24'h0000ff;
assign target7[156] = 24'h0000ff;
assign target7[157] = 24'h0000ff;
assign target7[158] = 24'h0000ff;
assign target7[159] = 24'h0000ff;
assign target7[160] = 24'h00ffff;
assign target7[161] = 24'h00ffff;
assign target7[162] = 24'h00ffff;
assign target7[163] = 24'h00ffff;
assign target7[164] = 24'h00ffff;
assign target7[165] = 24'h00ffff;
assign target7[166] = 24'h00ffff;
assign target7[167] = 24'h00ffff;
assign target7[168] = 24'h00ffff;
assign target7[169] = 24'h00ffff;
assign target7[170] = 24'h00ffff;
assign target7[171] = 24'h00ffff;
assign target7[172] = 24'h00ffff;
assign target7[173] = 24'h00ffff;
assign target7[174] = 24'h00ffff;
assign target7[175] = 24'h00ffff;
assign target7[176] = 24'h00ffff;
assign target7[177] = 24'h00ffff;
assign target7[178] = 24'h00ffff;
assign target7[179] = 24'h00ffff;
assign target7[180] = 24'hff00ff;
assign target7[181] = 24'hff00ff;
assign target7[182] = 24'hff00ff;
assign target7[183] = 24'hff00ff;
assign target7[184] = 24'hff00ff;
assign target7[185] = 24'hff00ff;
assign target7[186] = 24'hff00ff;
assign target7[187] = 24'hff00ff;
assign target7[188] = 24'hff00ff;
assign target7[189] = 24'hff00ff;
assign target7[190] = 24'hff00ff;
assign target7[191] = 24'hff00ff;
assign target7[192] = 24'hff00ff;
assign target7[193] = 24'hff00ff;
assign target7[194] = 24'hff00ff;
assign target7[195] = 24'hff00ff;
assign target7[196] = 24'hff00ff;
assign target7[197] = 24'hff00ff;
assign target7[198] = 24'hff00ff;
assign target7[199] = 24'hff00ff;
assign target7[200] = 24'hffff00;
assign target7[201] = 24'hffff00;
assign target7[202] = 24'hffff00;
assign target7[203] = 24'hffff00;
assign target7[204] = 24'hffff00;
assign target7[205] = 24'hffff00;
assign target7[206] = 24'hffff00;
assign target7[207] = 24'hffff00;
assign target7[208] = 24'hffff00;
assign target7[209] = 24'hffff00;
assign target7[210] = 24'hffff00;
assign target7[211] = 24'hffff00;
assign target7[212] = 24'hffff00;
assign target7[213] = 24'hffff00;
assign target7[214] = 24'hffff00;
assign target7[215] = 24'hffff00;
assign target7[216] = 24'hffff00;
assign target7[217] = 24'hffff00;
assign target7[218] = 24'hffff00;
assign target7[219] = 24'hffff00;
assign target7[220] = 24'h8f8f8f;
assign target7[221] = 24'h8f8f8f;
assign target7[222] = 24'h8f8f8f;
assign target7[223] = 24'h8f8f8f;
assign target7[224] = 24'h8f8f8f;
assign target7[225] = 24'h8f8f8f;
assign target7[226] = 24'h8f8f8f;
assign target7[227] = 24'h8f8f8f;
assign target7[228] = 24'h8f8f8f;
assign target7[229] = 24'h8f8f8f;
assign target7[230] = 24'h8f8f8f;
assign target7[231] = 24'h8f8f8f;
assign target7[232] = 24'h8f8f8f;
assign target7[233] = 24'h8f8f8f;
assign target7[234] = 24'h8f8f8f;
assign target7[235] = 24'h8f8f8f;
assign target7[236] = 24'h8f8f8f;
assign target7[237] = 24'h8f8f8f;
assign target7[238] = 24'h8f8f8f;
assign target7[239] = 24'h8f8f8f;
assign target7[240] = 24'h7a0000;
assign target7[241] = 24'h7a0000;
assign target7[242] = 24'h7a0000;
assign target7[243] = 24'h7a0000;
assign target7[244] = 24'h7a0000;
assign target7[245] = 24'h7a0000;
assign target7[246] = 24'h7a0000;
assign target7[247] = 24'h7a0000;
assign target7[248] = 24'h7a0000;
assign target7[249] = 24'h7a0000;
assign target7[250] = 24'h7a0000;
assign target7[251] = 24'h7a0000;
assign target7[252] = 24'h7a0000;
assign target7[253] = 24'h7a0000;
assign target7[254] = 24'h7a0000;
assign target7[255] = 24'h7a0000;
assign target7[256] = 24'h7a0000;
assign target7[257] = 24'h7a0000;
assign target7[258] = 24'h7a0000;
assign target7[259] = 24'h7a0000;
assign target7[260] = 24'h007a00;
assign target7[261] = 24'h007a00;
assign target7[262] = 24'h007a00;
assign target7[263] = 24'h007a00;
assign target7[264] = 24'h007a00;
assign target7[265] = 24'h007a00;
assign target7[266] = 24'h007a00;
assign target7[267] = 24'h007a00;
assign target7[268] = 24'h007a00;
assign target7[269] = 24'h007a00;
assign target7[270] = 24'h007a00;
assign target7[271] = 24'h007a00;
assign target7[272] = 24'h007a00;
assign target7[273] = 24'h007a00;
assign target7[274] = 24'h007a00;
assign target7[275] = 24'h007a00;
assign target7[276] = 24'h007a00;
assign target7[277] = 24'h007a00;
assign target7[278] = 24'h007a00;
assign target7[279] = 24'h007a00;
assign target7[280] = 24'h00008b;
assign target7[281] = 24'h00008b;
assign target7[282] = 24'h00008b;
assign target7[283] = 24'h00008b;
assign target7[284] = 24'h00008b;
assign target7[285] = 24'h00008b;
assign target7[286] = 24'h00008b;
assign target7[287] = 24'h00008b;
assign target7[288] = 24'h00008b;
assign target7[289] = 24'h00008b;
assign target7[290] = 24'h00008b;
assign target7[291] = 24'h00008b;
assign target7[292] = 24'h00008b;
assign target7[293] = 24'h00008b;
assign target7[294] = 24'h00008b;
assign target7[295] = 24'h00008b;
assign target7[296] = 24'h00008b;
assign target7[297] = 24'h00008b;
assign target7[298] = 24'h00008b;
assign target7[299] = 24'h00008b;
assign target7[300] = 24'h0088ff;
assign target7[301] = 24'h0088ff;
assign target7[302] = 24'h0088ff;
assign target7[303] = 24'h0088ff;
assign target7[304] = 24'h0088ff;
assign target7[305] = 24'h0088ff;
assign target7[306] = 24'h0088ff;
assign target7[307] = 24'h0088ff;
assign target7[308] = 24'h0088ff;
assign target7[309] = 24'h0088ff;
assign target7[310] = 24'h0088ff;
assign target7[311] = 24'h0088ff;
assign target7[312] = 24'h0088ff;
assign target7[313] = 24'h0088ff;
assign target7[314] = 24'h0088ff;
assign target7[315] = 24'h0088ff;
assign target7[316] = 24'h0088ff;
assign target7[317] = 24'h0088ff;
assign target7[318] = 24'h0088ff;
assign target7[319] = 24'h0088ff;
assign target7[320] = 24'h7100ff;
assign target7[321] = 24'h7100ff;
assign target7[322] = 24'h7100ff;
assign target7[323] = 24'h7100ff;
assign target7[324] = 24'h7100ff;
assign target7[325] = 24'h7100ff;
assign target7[326] = 24'h7100ff;
assign target7[327] = 24'h7100ff;
assign target7[328] = 24'h7100ff;
assign target7[329] = 24'h7100ff;
assign target7[330] = 24'h7100ff;
assign target7[331] = 24'h7100ff;
assign target7[332] = 24'h7100ff;
assign target7[333] = 24'h7100ff;
assign target7[334] = 24'h7100ff;
assign target7[335] = 24'h7100ff;
assign target7[336] = 24'h7100ff;
assign target7[337] = 24'h7100ff;
assign target7[338] = 24'h7100ff;
assign target7[339] = 24'h7100ff;
assign target7[340] = 24'h82ff00;
assign target7[341] = 24'h82ff00;
assign target7[342] = 24'h82ff00;
assign target7[343] = 24'h82ff00;
assign target7[344] = 24'h82ff00;
assign target7[345] = 24'h82ff00;
assign target7[346] = 24'h82ff00;
assign target7[347] = 24'h82ff00;
assign target7[348] = 24'h82ff00;
assign target7[349] = 24'h82ff00;
assign target7[350] = 24'h82ff00;
assign target7[351] = 24'h82ff00;
assign target7[352] = 24'h82ff00;
assign target7[353] = 24'h82ff00;
assign target7[354] = 24'h82ff00;
assign target7[355] = 24'h82ff00;
assign target7[356] = 24'h82ff00;
assign target7[357] = 24'h82ff00;
assign target7[358] = 24'h82ff00;
assign target7[359] = 24'h82ff00;
assign target7[360] = 24'h00ff74;
assign target7[361] = 24'h00ff74;
assign target7[362] = 24'h00ff74;
assign target7[363] = 24'h00ff74;
assign target7[364] = 24'h00ff74;
assign target7[365] = 24'h00ff74;
assign target7[366] = 24'h00ff74;
assign target7[367] = 24'h00ff74;
assign target7[368] = 24'h00ff74;
assign target7[369] = 24'h00ff74;
assign target7[370] = 24'h00ff74;
assign target7[371] = 24'h00ff74;
assign target7[372] = 24'h00ff74;
assign target7[373] = 24'h00ff74;
assign target7[374] = 24'h00ff74;
assign target7[375] = 24'h00ff74;
assign target7[376] = 24'h00ff74;
assign target7[377] = 24'h00ff74;
assign target7[378] = 24'h00ff74;
assign target7[379] = 24'h00ff74;
assign target7[380] = 24'hff007d;
assign target7[381] = 24'hff007d;
assign target7[382] = 24'hff007d;
assign target7[383] = 24'hff007d;
assign target7[384] = 24'hff007d;
assign target7[385] = 24'hff007d;
assign target7[386] = 24'hff007d;
assign target7[387] = 24'hff007d;
assign target7[388] = 24'hff007d;
assign target7[389] = 24'hff007d;
assign target7[390] = 24'hff007d;
assign target7[391] = 24'hff007d;
assign target7[392] = 24'hff007d;
assign target7[393] = 24'hff007d;
assign target7[394] = 24'hff007d;
assign target7[395] = 24'hff007d;
assign target7[396] = 24'hff007d;
assign target7[397] = 24'hff007d;
assign target7[398] = 24'hff007d;
assign target7[399] = 24'hff007d;
